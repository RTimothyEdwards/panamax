magic
tech sky130A
magscale 1 2
timestamp 1746115413
<< checkpaint >>
rect 39927 520724 40459 644952
rect 38963 519210 41531 520724
rect 38620 516642 41531 519210
rect 38620 515968 41188 516642
rect 38620 513400 41664 515968
rect 38904 512032 41664 513400
rect 38904 510244 41472 512032
rect 38904 507676 41644 510244
rect 39927 380104 40459 507676
<< metal2 >>
rect 40044 642702 40092 644952
rect 40044 609702 40092 611952
rect 40044 576702 40092 578952
rect 40044 541116 40092 545970
rect 40044 541068 40271 541116
rect 40223 519106 40271 541068
rect 39927 519058 40271 519106
rect 40223 517950 40271 519058
rect 39880 517902 40271 517950
rect 39880 514708 39928 517902
rect 39880 514660 40404 514708
rect 40356 513340 40404 514660
rect 40164 513292 40404 513340
rect 40164 508984 40212 513292
rect 40164 508936 40459 508984
rect 40411 481036 40459 508936
rect 40044 480988 40459 481036
rect 40044 479120 40092 480988
rect 40044 446104 40092 448356
rect 40044 413104 40092 415356
rect 40044 380104 40092 382356
<< properties >>
string flatten true
<< end >>
