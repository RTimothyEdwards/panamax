magic
tech sky130A
magscale 1 2
timestamp 1746202612
<< metal4 >>
rect 142 140 16102 560
<< metal5 >>
rect 9102 15260 9452 15400
tri 8192 15120 8332 15260 se
rect 8332 15120 9452 15260
tri 8052 14840 8192 14980 se
rect 8192 14840 9452 15120
tri 6892 14700 7032 14840 se
rect 7032 14700 8542 14840
rect 6892 14630 8542 14700
tri 6752 14420 6892 14560 se
rect 6892 14490 8402 14630
tri 8402 14490 8542 14630 nw
rect 6892 14420 7212 14490
tri 7212 14420 7282 14490 nw
rect 6302 14210 7212 14420
rect 9102 14350 9452 14840
rect 9102 14280 10922 14350
rect 6302 14070 7072 14210
tri 7072 14070 7212 14210 nw
tri 8542 14140 8682 14280 se
rect 8682 14140 10922 14280
tri 7772 14070 7842 14140 se
rect 7842 14070 10922 14140
tri 7142 13440 7772 14070 se
rect 7772 14000 10922 14070
rect 7772 13580 10642 14000
tri 10642 13860 10782 14000 nw
rect 7772 13440 10502 13580
tri 10502 13440 10642 13580 nw
tri 7002 12880 7142 13020 se
rect 7142 12880 10502 13440
rect 7002 12600 10502 12880
tri 10502 12600 10642 12740 sw
rect 4062 11620 4412 12320
rect 7002 12040 10642 12600
tri 7002 11900 7142 12040 ne
rect 7142 11900 10642 12040
tri 10642 11900 10922 12180 sw
rect 7142 11760 8542 11900
tri 8542 11760 8682 11900 nw
rect 9102 11760 10922 11900
rect 7142 11620 7975 11760
rect 3642 11200 4762 11620
tri 3642 11060 3782 11200 ne
rect 3782 10780 4622 11200
tri 4622 11060 4762 11200 nw
tri 7142 11107 7655 11620 ne
rect 7655 11107 7975 11620
tri 7975 11543 8192 11760 nw
rect 9102 10990 9522 11760
tri 10222 11480 10502 11760 ne
rect 10502 11480 10922 11760
tri 14842 11620 15262 12040 se
rect 15262 11620 15582 12040
tri 14702 11480 14842 11620 se
tri 14422 11200 14702 11480 se
rect 14702 11200 14842 11480
tri 14212 10990 14422 11200 se
rect 14422 10990 14842 11200
tri 14842 11060 15402 11620 nw
rect 9102 10920 11902 10990
tri 8542 10780 8682 10920 se
rect 8682 10780 11902 10920
rect 4062 10430 4412 10780
rect 7422 10640 11902 10780
tri 13862 10640 14212 10990 se
rect 14212 10920 14842 10990
rect 14212 10640 14702 10920
tri 14702 10780 14842 10920 nw
tri 7352 10430 7422 10500 se
rect 7422 10430 11202 10640
rect 4062 10360 5602 10430
tri 7282 10360 7352 10430 se
rect 7352 10360 11202 10430
tri 11202 10360 11482 10640 nw
tri 13722 10500 13862 10640 se
rect 13862 10500 14702 10640
tri 2942 10220 3082 10360 se
rect 3082 10220 5602 10360
rect 2102 10080 5602 10220
tri 6862 10080 7142 10360 se
rect 7142 10080 11202 10360
tri 1402 9240 2102 9940 se
rect 2102 9380 5042 10080
tri 5042 9940 5182 10080 nw
tri 6722 9940 6862 10080 se
rect 6862 9940 10782 10080
rect 2102 9240 4902 9380
tri 4902 9240 5042 9380 nw
tri 6022 9240 6722 9940 se
rect 6722 9240 10782 9940
tri 10782 9660 11202 10080 nw
rect 12672 10010 13022 10500
tri 13442 10220 13722 10500 se
rect 13722 10220 14562 10500
tri 14562 10360 14702 10500 nw
tri 13372 10010 13442 10080 se
rect 13442 10010 14562 10220
rect 12672 9800 14562 10010
tri 1262 8680 1402 8820 se
rect 1402 8680 4902 9240
rect 1262 8120 4902 8680
tri 5462 8540 6022 9100 se
rect 6022 8540 10642 9240
tri 10642 9100 10782 9240 nw
tri 12532 9240 12672 9380 se
rect 12672 9240 14422 9800
tri 14422 9660 14562 9800 nw
tri 12462 9100 12532 9170 se
rect 12532 9100 14422 9240
tri 4902 8120 5042 8260 sw
rect 1262 7420 5042 8120
tri 1262 7280 1402 7420 ne
rect 1402 6860 5042 7420
tri 1402 6650 1612 6860 ne
rect 1612 6720 5042 6860
tri 5392 7910 5462 7980 se
rect 5462 7910 10642 8540
rect 5392 6860 10642 7910
tri 11622 8120 12462 8960 se
rect 12462 8120 14282 9100
tri 14282 8960 14422 9100 nw
tri 11342 7560 11622 7840 se
rect 11622 7560 14282 8120
tri 11132 7280 11342 7490 se
rect 11342 7280 14282 7560
tri 10992 6860 11132 7000 se
rect 11132 6860 14282 7280
rect 5392 6720 14282 6860
tri 14282 6720 14422 6860 sw
rect 1612 6650 3082 6720
rect 282 6580 702 6650
tri 702 6580 772 6650 sw
tri 1612 6580 1682 6650 ne
rect 1682 6580 3082 6650
tri 3082 6580 3222 6720 nw
tri 3642 6580 3782 6720 ne
rect 3782 6580 14422 6720
rect 282 6440 842 6580
tri 842 6440 982 6580 sw
tri 1682 6440 1822 6580 ne
rect 1822 6440 2662 6580
rect 282 6300 1122 6440
tri 562 6120 742 6300 ne
rect 742 6160 1122 6300
tri 1122 6160 1402 6440 sw
rect 1962 6160 2662 6440
tri 2662 6300 2942 6580 nw
rect 4062 6440 14422 6580
rect 742 6120 1542 6160
tri 882 5840 1162 6120 ne
rect 1162 6090 1542 6120
tri 1542 6090 1612 6160 sw
rect 1962 6090 2592 6160
tri 2592 6090 2662 6160 nw
rect 1162 5840 2592 6090
tri 1302 5740 1402 5840 ne
rect 1402 5740 2592 5840
tri 1542 5600 1682 5740 ne
rect 1682 5600 3422 5740
tri 1822 5460 1962 5600 ne
rect 1962 5460 3422 5600
tri 3422 5460 3702 5740 sw
rect 4062 5460 4482 6440
tri 4842 6300 4982 6440 ne
rect 4982 6300 14422 6440
tri 5042 6020 5322 6300 ne
rect 5322 6020 14422 6300
rect 1962 5180 4482 5460
rect 5322 5880 11762 6020
tri 11762 5880 11902 6020 nw
rect 5322 5740 11342 5880
tri 11342 5740 11482 5880 nw
tri 5322 5180 5882 5740 ne
rect 5882 5220 11342 5740
tri 11342 5220 11622 5500 sw
rect 5882 5180 11622 5220
rect 2242 5040 4482 5180
tri 4482 5040 4622 5180 sw
rect 5882 5040 8402 5180
tri 8402 5040 8542 5180 nw
tri 8962 5040 9102 5180 ne
rect 9102 5040 11622 5180
tri 2242 4900 2382 5040 ne
rect 2382 4900 4902 5040
tri 4902 4900 5042 5040 sw
tri 2662 4060 3502 4900 ne
rect 3502 3780 5462 4900
rect 5882 4760 7282 5040
tri 7282 4900 7422 5040 nw
tri 5882 4340 6302 4760 ne
rect 6302 4340 6862 4760
tri 6862 4340 7282 4760 nw
rect 9242 4760 11622 5040
tri 5462 3780 6022 4340 sw
tri 6302 4200 6442 4340 ne
rect 6442 3780 6862 4340
tri 3362 3500 3502 3640 se
rect 3502 3500 6862 3780
rect 3362 3360 6862 3500
tri 6862 3360 7282 3780 sw
rect 3362 3220 7562 3360
tri 7562 3220 7702 3360 sw
rect 3362 3080 8122 3220
tri 8122 3080 8262 3220 sw
rect 9242 3080 9802 4760
tri 10222 4620 10362 4760 ne
rect 10362 4620 11622 4760
tri 11622 4620 12042 5040 sw
tri 10922 4340 11202 4620 ne
rect 11202 4480 12042 4620
rect 12602 4480 13022 6020
tri 13442 5880 13582 6020 ne
rect 13582 5880 14422 6020
tri 14422 5880 14702 6160 sw
tri 13822 5320 14382 5880 ne
rect 14382 5320 14702 5880
tri 13722 4620 14002 4900 se
rect 14002 4760 15262 4900
tri 15262 4760 15402 4900 sw
rect 14002 4620 15402 4760
tri 13442 4480 13582 4620 se
rect 13582 4480 15402 4620
rect 11202 4410 15402 4480
rect 11202 4340 15262 4410
tri 11622 4060 11902 4340 ne
rect 11902 4060 15262 4340
rect 11902 3710 16102 4060
rect 11902 3640 15402 3710
tri 10922 3080 11482 3640 se
rect 11482 3500 15402 3640
rect 11482 3080 15262 3500
tri 15262 3360 15402 3500 nw
rect 3362 2800 15262 3080
rect 3362 2660 7212 2800
tri 3362 2520 3502 2660 ne
rect 3502 2380 7212 2660
rect 7562 2660 15262 2800
rect 7562 2380 8052 2660
rect 3502 2240 8052 2380
rect 8402 2520 14982 2660
tri 14982 2520 15122 2660 nw
rect 8402 2240 8962 2520
rect 3502 2100 8962 2240
rect 9312 2100 9802 2520
rect 10152 2100 10642 2520
rect 10992 2100 14982 2520
rect 3502 1960 14982 2100
tri 3502 1820 3642 1960 ne
rect 3642 1540 14842 1960
tri 14842 1820 14982 1960 nw
tri 3642 1400 3782 1540 ne
rect 3782 1260 14422 1540
tri 3782 840 4202 1260 ne
rect 4202 700 14422 1260
tri 14422 1120 14842 1540 nw
tri 4202 560 4342 700 ne
rect 4342 560 14422 700
<< fillblock >>
rect 2 10360 16262 15560
rect 0 9800 16262 10360
rect 2 0 16262 9800
<< end >>
