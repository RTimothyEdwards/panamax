magic
tech sky130A
magscale 1 2
timestamp 1726839386
<< checkpaint >>
rect -335 -3690 3913 1114
<< metal1 >>
rect 753 4232 759 4444
rect 811 4284 817 4444
rect 811 4232 893 4284
<< via1 >>
rect 759 4232 811 4444
<< metal2 >>
rect 270 9992 318 16814
rect 266 9983 322 9992
rect 266 9825 322 9835
rect 270 -2001 318 9825
rect 364 -1467 412 16814
rect 458 -1014 510 16814
rect 556 481 604 16814
rect 545 461 617 481
rect 545 381 617 401
rect 448 -1037 520 -1014
rect 448 -1119 520 -1097
rect 349 -1487 421 -1467
rect 349 -1572 421 -1547
rect 364 -2001 412 -1572
rect 458 -2001 510 -1119
rect 556 -2001 604 381
rect 652 183 700 16814
rect 774 16259 834 16268
rect 834 16049 845 16095
rect 774 16030 834 16039
rect 774 15856 834 15865
rect 834 15640 845 15686
rect 774 15627 834 15636
rect 745 15535 845 15544
rect 805 15492 845 15535
rect 745 15306 805 15315
rect 765 14379 835 14384
rect 761 14159 770 14379
rect 830 14219 840 14379
rect 830 14167 843 14219
rect 830 14159 839 14167
rect 765 14154 835 14159
rect 755 13659 825 13664
rect 751 13439 760 13659
rect 820 13508 830 13659
rect 820 13456 842 13508
rect 820 13447 830 13456
rect 820 13439 829 13447
rect 755 13434 825 13439
rect 765 12549 835 12554
rect 761 12329 770 12549
rect 830 12329 840 12549
rect 761 12299 840 12329
rect 761 12247 862 12299
rect 737 11390 746 11610
rect 806 11450 815 11610
rect 806 11398 853 11450
rect 806 11390 815 11398
rect 773 10938 782 11158
rect 842 11072 851 11158
rect 842 11020 868 11072
rect 842 10938 851 11020
rect 767 10786 827 10795
rect 827 10568 868 10620
rect 767 10557 827 10566
rect 761 10409 821 10419
rect 821 10355 842 10407
rect 761 10180 821 10189
rect 763 9794 833 9803
rect 763 9574 768 9794
rect 828 9678 833 9794
rect 828 9626 842 9678
rect 828 9574 833 9626
rect 763 9565 833 9574
rect 770 9343 830 9347
rect 765 9338 835 9343
rect 765 9118 770 9338
rect 830 9118 835 9338
rect 765 9092 835 9118
rect 765 9040 842 9092
rect 758 7665 767 7885
rect 827 7721 836 7885
rect 827 7669 851 7721
rect 827 7665 836 7669
rect 769 7045 839 7054
rect 769 6825 774 7045
rect 834 6825 839 7045
rect 769 6799 839 6825
rect 769 6747 844 6799
rect 755 4835 815 4844
rect 755 4606 815 4615
rect 759 4444 811 4606
rect 759 4226 811 4232
rect 760 3347 769 3567
rect 829 3403 838 3567
rect 829 3351 859 3403
rect 829 3347 838 3351
rect 758 2825 767 3113
rect 855 2825 865 3113
rect 768 1419 777 1707
rect 865 1419 875 1707
rect 768 1386 875 1419
rect 794 1250 1050 1259
rect 1014 1190 1050 1250
rect 794 1181 1050 1190
rect 756 989 842 1029
rect 756 555 796 989
rect 741 546 801 555
rect 741 317 801 326
rect 892 322 932 827
rect 641 163 713 183
rect 641 82 713 103
rect 866 102 875 322
rect 935 102 944 322
rect 652 -2001 700 82
<< via2 >>
rect 266 9835 322 9983
rect 545 401 617 461
rect 448 -1097 520 -1037
rect 349 -1547 421 -1487
rect 774 16039 834 16259
rect 774 15636 834 15856
rect 745 15315 805 15535
rect 770 14159 830 14379
rect 760 13439 820 13659
rect 770 12329 830 12549
rect 746 11390 806 11610
rect 782 10938 842 11158
rect 767 10566 827 10786
rect 761 10189 821 10409
rect 768 9574 828 9794
rect 770 9118 830 9338
rect 767 7665 827 7885
rect 774 6825 834 7045
rect 755 4615 815 4835
rect 769 3347 829 3567
rect 767 2825 855 3113
rect 777 1419 865 1707
rect 794 1190 1014 1250
rect 741 326 801 546
rect 641 103 713 163
rect 875 102 935 322
<< metal3 >>
rect 0 16566 842 16690
rect 769 16259 839 16275
rect 769 16108 774 16259
rect 0 16039 774 16108
rect 834 16039 839 16259
rect 0 16038 839 16039
rect 769 16034 839 16038
rect 769 15856 839 15871
rect 769 15698 774 15856
rect 0 15636 774 15698
rect 834 15636 839 15856
rect 0 15628 839 15636
rect 458 15535 810 15554
rect 458 15484 745 15535
rect 458 15354 528 15484
rect 0 15284 528 15354
rect 740 15315 745 15484
rect 805 15315 810 15535
rect 740 15310 810 15315
rect 0 14422 835 14492
rect 765 14379 835 14422
rect 765 14159 770 14379
rect 830 14159 835 14379
rect 765 14154 835 14159
rect 0 13702 825 13772
rect 755 13659 825 13702
rect 755 13439 760 13659
rect 820 13439 825 13659
rect 755 13434 825 13439
rect 0 12549 835 12572
rect 0 12502 770 12549
rect 765 12329 770 12502
rect 830 12329 835 12549
rect 765 12324 835 12329
rect 0 11730 811 11800
rect 741 11610 811 11730
rect 741 11390 746 11610
rect 806 11390 811 11610
rect 741 11385 811 11390
rect 0 11246 564 11316
rect 494 11162 564 11246
rect 777 11162 847 11163
rect 494 11158 847 11162
rect 494 11092 782 11158
rect 777 10938 782 11092
rect 842 10938 847 11158
rect 777 10933 847 10938
rect 0 10802 832 10872
rect 762 10786 832 10802
rect 762 10566 767 10786
rect 827 10566 832 10786
rect 762 10560 832 10566
rect 756 10409 826 10414
rect 756 10254 761 10409
rect 0 10189 761 10254
rect 821 10189 826 10409
rect 0 10184 826 10189
rect 261 9983 327 9992
rect 261 9835 266 9983
rect 322 9835 327 9983
rect 261 9800 327 9835
rect 0 9794 833 9800
rect 0 9730 768 9794
rect 763 9574 768 9730
rect 828 9574 833 9794
rect 763 9569 833 9574
rect 0 9343 770 9344
rect 0 9338 835 9343
rect 0 9274 770 9338
rect 765 9118 770 9274
rect 830 9118 835 9338
rect 765 9113 835 9118
rect 0 8108 827 8178
rect 767 7890 827 8108
rect 762 7885 832 7890
rect 762 7665 767 7885
rect 827 7665 832 7885
rect 762 7660 832 7665
rect 0 7528 851 7598
rect 0 7045 839 7050
rect 0 6980 774 7045
rect 769 6825 774 6980
rect 834 6825 839 7045
rect 769 6820 839 6825
rect 750 4838 820 4840
rect 0 4835 820 4838
rect 0 4768 755 4835
rect 750 4615 755 4768
rect 815 4615 820 4835
rect 750 4610 820 4615
rect 0 3992 842 4206
rect 0 3572 834 3642
rect 764 3567 834 3572
rect 764 3347 769 3567
rect 829 3347 834 3567
rect 764 3342 834 3347
rect 762 3113 860 3118
rect 762 3112 767 3113
rect 0 2982 767 3112
rect 762 2825 767 2982
rect 855 2825 860 3113
rect 762 2820 860 2825
rect 772 1707 870 1713
rect 772 1680 777 1707
rect 0 1552 777 1680
rect 772 1419 777 1552
rect 865 1419 870 1707
rect 772 1414 870 1419
rect 0 1262 846 1332
rect 776 1255 846 1262
rect 776 1250 1074 1255
rect 776 1190 794 1250
rect 1014 1190 1074 1250
rect 776 1185 1074 1190
rect 0 988 842 1058
rect 657 852 1005 922
rect 657 746 727 852
rect 4 676 727 746
rect 736 546 806 556
rect 736 466 741 546
rect 0 461 741 466
rect 0 401 545 461
rect 617 401 741 461
rect 0 396 741 401
rect 736 326 741 396
rect 801 326 806 546
rect 736 321 806 326
rect 870 322 940 327
rect 870 168 875 322
rect 0 163 875 168
rect 0 103 641 163
rect 713 103 875 163
rect 0 102 875 103
rect 935 102 940 322
rect 0 98 940 102
rect 870 97 940 98
rect 2653 -212 3552 -202
rect 2653 -374 2657 -212
rect 3540 -374 3552 -212
rect 2653 -382 3552 -374
rect 2653 -710 10095 -702
rect 2653 -876 9167 -710
rect 10079 -876 10095 -710
rect 2653 -882 10095 -876
rect 0 -1037 942 -1032
rect 0 -1097 448 -1037
rect 520 -1097 942 -1037
rect 0 -1102 942 -1097
rect 2653 -1209 3552 -1202
rect 2653 -1371 2657 -1209
rect 3540 -1371 3552 -1209
rect 2653 -1382 3552 -1371
rect 0 -1487 952 -1482
rect 0 -1547 349 -1487
rect 421 -1547 952 -1487
rect 0 -1552 952 -1547
rect 2653 -1709 10095 -1702
rect 2653 -1875 9167 -1709
rect 10079 -1875 10095 -1709
rect 2653 -1882 10095 -1875
rect 2653 -2209 3552 -2202
rect 2653 -2371 2656 -2209
rect 3539 -2371 3552 -2209
rect 2653 -2382 3552 -2371
<< via3 >>
rect 2657 -374 3540 -212
rect 9167 -876 10079 -710
rect 2657 -1371 3540 -1209
rect 9167 -1875 10079 -1709
rect 2656 -2371 3539 -2209
<< metal4 >>
rect 2655 -212 3542 -210
rect 2655 -374 2657 -212
rect 3540 -374 3542 -212
rect 2655 -376 3542 -374
rect 9165 -710 10081 -708
rect 9165 -876 9167 -710
rect 10079 -876 10081 -710
rect 9165 -878 10081 -876
rect 2655 -1209 3542 -1207
rect 2655 -1371 2657 -1209
rect 3540 -1371 3542 -1209
rect 2655 -1373 3542 -1371
rect 9165 -1709 10081 -1707
rect 9165 -1875 9167 -1709
rect 10079 -1875 10081 -1709
rect 9165 -1877 10081 -1875
rect 2654 -2209 3541 -2207
rect 2654 -2371 2656 -2209
rect 3539 -2371 3541 -2209
rect 2654 -2373 3541 -2371
use constant_block  constant_block_0
timestamp 1706127523
transform 0 -1 3149 -1 0 0
box 146 496 2430 2224
<< labels >>
flabel metal3 s 0 98 300 168 0 FreeSans 320 0 0 0 tie_lo_esd
port 1 nsew
flabel metal3 s 0 988 300 1058 0 FreeSans 320 0 0 0 enable_vddio
port 4 nsew
flabel metal3 s 0 1262 300 1332 0 FreeSans 320 0 0 0 slow
port 5 nsew
flabel metal3 s 0 1552 300 1680 0 FreeSans 320 0 0 0 pad_a_esd_0_h
port 6 nsew
flabel metal3 s 0 2982 300 3112 0 FreeSans 320 0 0 0 pad_a_esd_1_h
port 7 nsew
flabel metal3 s 0 3572 300 3642 0 FreeSans 320 0 0 0 dm[1]
port 8 nsew
flabel metal3 s 0 3992 300 4206 0 FreeSans 320 0 0 0 pad_a_noesd_h
port 9 nsew
flabel metal3 s 0 4768 300 4838 0 FreeSans 320 0 0 0 analog_en
port 10 nsew
flabel metal3 s 0 6980 300 7050 0 FreeSans 320 0 0 0 dm[0]
port 11 nsew
flabel metal3 s 0 7528 300 7598 0 FreeSans 320 0 0 0 analog_pol
port 12 nsew
flabel metal3 s 0 8108 300 8178 0 FreeSans 320 0 0 0 inp_dis
port 13 nsew
flabel metal3 s 0 9274 300 9344 0 FreeSans 320 0 0 0 enable_inp_h
port 14 nsew
flabel metal3 s 0 9730 300 9800 0 FreeSans 320 0 0 0 enable_h
port 15 nsew
flabel metal3 s 0 10184 300 10254 0 FreeSans 320 0 0 0 hld_h_n
port 16 nsew
flabel metal3 s 0 10802 300 10872 0 FreeSans 320 0 0 0 analog_sel
port 17 nsew
flabel metal3 s 0 11246 300 11316 0 FreeSans 320 0 0 0 dm[2]
port 18 nsew
flabel metal3 s 0 11730 300 11800 0 FreeSans 320 0 0 0 hld_ovr
port 19 nsew
flabel metal3 s 0 12502 300 12572 0 FreeSans 320 0 0 0 out
port 20 nsew
flabel metal3 s 0 13702 300 13772 0 FreeSans 320 0 0 0 enable_vswitch_h
port 21 nsew
flabel metal3 s 0 14422 300 14492 0 FreeSans 320 0 0 0 enable_vdda_h
port 22 nsew
flabel metal3 s 0 15628 300 15698 0 FreeSans 320 0 0 0 ib_mode_sel
port 24 nsew
flabel metal3 s 0 16038 300 16108 0 FreeSans 320 0 0 0 oe_n
port 25 nsew
flabel metal3 s 0 16566 300 16690 0 FreeSans 320 0 0 0 in_h
port 26 nsew
flabel metal3 s 0 -1552 300 -1482 0 FreeSans 320 0 0 0 one
port 27 nsew
flabel metal3 s 0 -1102 300 -1032 0 FreeSans 320 0 0 0 zero
port 28 nsew
flabel metal3 s 0 15284 300 15354 0 FreeSans 320 0 0 0 vtrip_sel
port 23 nsew
flabel metal3 s 0 396 300 466 0 FreeSans 320 0 0 0 tie_hi_esd
port 3 nsew
flabel metal3 s 4 676 304 746 0 FreeSans 320 0 0 0 in
port 2 nsew
<< properties >>
string FIXED_BBOX 0 770 1249 16770
string flatten true
<< end >>
