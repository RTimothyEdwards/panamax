magic
tech sky130A
magscale 1 2
timestamp 1746117482
<< checkpaint >>
rect 2024 4996 4600 5060
rect 2024 4834 5748 4996
rect -1177 4774 5748 4834
rect -1570 -784 5748 4774
rect -1570 -898 5448 -784
rect -1366 -1318 5448 -898
rect -828 -1764 1978 -1318
<< isosubstrate >>
rect 260 560 3666 3400
<< viali >>
rect 1663 2610 1697 2644
rect 1951 2610 1985 2644
rect 2431 1944 2465 1978
<< metal1 >>
rect 480 3282 3456 3307
rect 480 3230 2122 3282
rect 2174 3230 2186 3282
rect 2238 3230 3456 3282
rect 480 3205 3456 3230
rect 1651 2644 1709 2650
rect 1651 2610 1663 2644
rect 1697 2641 1709 2644
rect 1939 2644 1997 2650
rect 1939 2641 1951 2644
rect 1697 2613 1951 2641
rect 1697 2610 1709 2613
rect 1651 2604 1709 2610
rect 1939 2610 1951 2613
rect 1985 2641 1997 2644
rect 3282 2641 3288 2653
rect 1985 2613 3288 2641
rect 1985 2610 1997 2613
rect 1939 2604 1997 2610
rect 3282 2601 3288 2613
rect 3340 2601 3346 2653
rect 480 2468 3456 2493
rect 480 2416 822 2468
rect 874 2416 886 2468
rect 938 2416 3456 2468
rect 480 2391 3456 2416
rect 1536 2286 2110 2289
rect 1536 2232 1670 2286
rect 1664 2226 1670 2232
rect 1854 2232 2110 2286
rect 1854 2226 1860 2232
rect 1664 2222 1860 2226
rect 592 1935 598 1987
rect 650 1975 656 1987
rect 2419 1978 2477 1984
rect 2419 1975 2431 1978
rect 650 1947 2431 1975
rect 650 1935 656 1947
rect 2419 1944 2431 1947
rect 2465 1944 2477 1978
rect 2419 1938 2477 1944
rect 480 1654 3456 1679
rect 480 1602 2122 1654
rect 2174 1602 2186 1654
rect 2238 1602 3456 1654
rect 480 1577 3456 1602
rect 480 840 3456 865
rect 480 788 822 840
rect 874 788 886 840
rect 938 788 3456 840
rect 480 763 3456 788
<< via1 >>
rect 2122 3230 2174 3282
rect 2186 3230 2238 3282
rect 3288 2601 3340 2653
rect 822 2416 874 2468
rect 886 2416 938 2468
rect 1670 2226 1854 2286
rect 598 1935 650 1987
rect 2122 1602 2174 1654
rect 2186 1602 2238 1654
rect 822 788 874 840
rect 886 788 938 840
<< metal2 >>
rect 2112 3284 2248 3307
rect 2168 3282 2192 3284
rect 2174 3230 2186 3282
rect 2168 3228 2192 3230
rect 2112 3205 2248 3228
rect 3288 2653 3340 2659
rect 3288 2595 3340 2601
rect 812 2470 948 2493
rect 868 2468 892 2470
rect 874 2416 886 2468
rect 868 2414 892 2416
rect 812 2391 948 2414
rect 1660 2286 1864 2296
rect 1660 2226 1670 2286
rect 1854 2226 1864 2286
rect 1660 2214 1864 2226
rect 598 1987 650 1993
rect 598 1929 650 1935
rect 610 800 638 1929
rect 2112 1656 2248 1679
rect 2168 1654 2192 1656
rect 2174 1602 2186 1654
rect 2168 1600 2192 1602
rect 2112 1577 2248 1600
rect 812 842 948 865
rect 868 840 892 842
rect 596 544 652 800
rect 874 788 886 840
rect 3301 800 3329 2595
rect 868 786 892 788
rect 812 763 948 786
rect 3288 544 3344 800
<< via2 >>
rect 2112 3282 2168 3284
rect 2192 3282 2248 3284
rect 2112 3230 2122 3282
rect 2122 3230 2168 3282
rect 2192 3230 2238 3282
rect 2238 3230 2248 3282
rect 2112 3228 2168 3230
rect 2192 3228 2248 3230
rect 812 2468 868 2470
rect 892 2468 948 2470
rect 812 2416 822 2468
rect 822 2416 868 2468
rect 892 2416 938 2468
rect 938 2416 948 2468
rect 812 2414 868 2416
rect 892 2414 948 2416
rect 1670 2226 1854 2286
rect 2112 1654 2168 1656
rect 2192 1654 2248 1656
rect 2112 1602 2122 1654
rect 2122 1602 2168 1654
rect 2192 1602 2238 1654
rect 2238 1602 2248 1654
rect 2112 1600 2168 1602
rect 2192 1600 2248 1602
rect 812 840 868 842
rect 892 840 948 842
rect 812 788 822 840
rect 822 788 868 840
rect 892 788 938 840
rect 938 788 948 840
rect 812 786 868 788
rect 892 786 948 788
<< metal3 >>
rect 790 2470 970 3307
rect 2090 3284 2270 3307
rect 790 2414 812 2470
rect 868 2414 892 2470
rect 948 2414 970 2470
rect 790 842 970 2414
rect 1670 2296 1850 3256
rect 2090 3228 2112 3284
rect 2168 3228 2192 3284
rect 2248 3228 2270 3284
rect 1660 2286 1864 2296
rect 1660 2226 1670 2286
rect 1854 2226 1864 2286
rect 1660 2214 1864 2226
rect 790 786 812 842
rect 868 786 892 842
rect 948 786 970 842
rect 1670 814 1850 2214
rect 2090 1656 2270 3228
rect 2090 1600 2112 1656
rect 2168 1600 2192 1656
rect 2248 1600 2270 1656
rect 790 763 970 786
rect 2090 763 2270 1600
rect 2970 814 3150 3256
use sky130_fd_sc_hvl__diode_2  ANTENNA_lvlshiftdown_A $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1738263620
transform 1 0 1536 0 -1 3256
box -66 -43 258 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1738263620
transform 1 0 480 0 -1 1628
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_8
timestamp 1738263620
transform 1 0 1248 0 -1 1628
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  FILLER_0_16
timestamp 1738263620
transform 1 0 2016 0 -1 1628
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1738263620
transform 1 0 2784 0 -1 1628
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_2  FILLER_0_28 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1738263620
transform 1 0 3168 0 -1 1628
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_1  FILLER_0_30 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1738263620
transform 1 0 3360 0 -1 1628
box -66 -43 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_1_0
timestamp 1738263620
transform 1 0 480 0 1 1628
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_4  FILLER_1_8
timestamp 1738263620
transform 1 0 1248 0 1 1628
box -66 -43 450 897
use sky130_fd_sc_hvl__fill_1  FILLER_1_12
timestamp 1738263620
transform 1 0 1632 0 1 1628
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  FILLER_1_30
timestamp 1738263620
transform 1 0 3360 0 1 1628
box -66 -43 162 897
use sky130_fd_sc_hvl__decap_8  FILLER_2_0
timestamp 1738263620
transform 1 0 480 0 -1 3256
box -66 -43 834 897
use sky130_fd_sc_hvl__fill_2  FILLER_2_8
timestamp 1738263620
transform 1 0 1248 0 -1 3256
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_1  FILLER_2_10
timestamp 1738263620
transform 1 0 1440 0 -1 3256
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_1  FILLER_2_30
timestamp 1738263620
transform 1 0 3360 0 -1 3256
box -66 -43 162 897
use sky130_fd_sc_hvl__lsbufhv2lv_1  lvlshiftdown $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1738263620
transform 1 0 1826 0 1 1628
box -66 -43 1698 1671
<< labels >>
flabel metal2 s 3288 544 3344 800 0 FreeSans 480 0 0 0 A
port 0 nsew signal input
flabel metal2 s 596 544 652 800 0 FreeSans 480 0 0 0 X
port 1 nsew signal tristate
flabel metal3 s 790 763 970 3307 0 FreeSans 640 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal3 s 2090 763 2270 3307 0 FreeSans 640 90 0 0 VGND
port 3 nsew ground bidirectional
flabel metal3 s 1670 814 1850 3256 0 FreeSans 640 90 0 0 LVPWR
port 4 nsew power bidirectional
flabel metal3 s 2970 814 3150 3256 0 FreeSans 640 90 0 0 LVGND
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 4000 3400
<< end >>
