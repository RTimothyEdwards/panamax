magic
tech sky130A
magscale 1 2
timestamp 1706127523
<< checkpaint >>
rect -1114 -764 3690 3484
<< viali >>
rect 899 1941 933 1975
rect 1067 1941 1101 1975
rect 1235 1941 1269 1975
rect 1403 1941 1437 1975
rect 1571 1941 1605 1975
rect 1739 1941 1773 1975
rect 1907 1941 1941 1975
rect 2075 1941 2109 1975
rect 2243 1941 2277 1975
rect 581 1853 615 1887
rect 899 1763 933 1797
rect 1067 1763 1101 1797
rect 1235 1763 1269 1797
rect 1403 1763 1437 1797
rect 1571 1763 1605 1797
rect 1739 1763 1773 1797
rect 1907 1763 1941 1797
rect 2075 1763 2109 1797
rect 2243 1763 2277 1797
rect 765 1513 799 1547
rect 581 1173 615 1207
rect 899 853 933 887
rect 1067 853 1101 887
rect 1235 853 1269 887
rect 1403 853 1437 887
rect 1571 853 1605 887
rect 1739 853 1773 887
rect 1907 853 1941 887
rect 2075 853 2109 887
rect 2243 853 2277 887
rect 581 765 615 799
rect 899 675 933 709
rect 1067 675 1101 709
rect 1235 675 1269 709
rect 1403 675 1437 709
rect 1571 675 1605 709
rect 1739 675 1773 709
rect 1907 675 1941 709
rect 2075 675 2109 709
rect 2243 675 2277 709
<< metal1 >>
rect 201 2202 2382 2224
rect 201 2150 234 2202
rect 286 2150 298 2202
rect 350 2150 1234 2202
rect 1286 2150 1298 2202
rect 1350 2150 2234 2202
rect 2286 2150 2298 2202
rect 2350 2150 2382 2202
rect 201 2128 2382 2150
rect 887 1975 2289 1981
rect 887 1941 899 1975
rect 933 1941 1067 1975
rect 1101 1941 1235 1975
rect 1269 1941 1403 1975
rect 1437 1941 1571 1975
rect 1605 1941 1739 1975
rect 1773 1941 1907 1975
rect 1941 1941 2075 1975
rect 2109 1941 2243 1975
rect 2277 1941 2289 1975
rect 887 1940 2289 1941
rect 887 1935 1400 1940
rect 566 1884 572 1896
rect 527 1856 572 1884
rect 566 1844 572 1856
rect 624 1844 630 1896
rect 1394 1803 1400 1935
rect 887 1797 1400 1803
rect 1452 1935 2289 1940
rect 1452 1803 1458 1935
rect 1452 1797 2289 1803
rect 887 1763 899 1797
rect 933 1763 1067 1797
rect 1101 1763 1235 1797
rect 1269 1768 1400 1797
rect 1452 1768 1571 1797
rect 1269 1763 1403 1768
rect 1437 1763 1571 1768
rect 1605 1763 1739 1797
rect 1773 1763 1907 1797
rect 1941 1763 2075 1797
rect 2109 1763 2243 1797
rect 2277 1763 2289 1797
rect 887 1757 2289 1763
rect 201 1658 2382 1680
rect 201 1606 734 1658
rect 786 1606 798 1658
rect 850 1606 1734 1658
rect 1786 1606 1798 1658
rect 1850 1606 2382 1658
rect 201 1584 2382 1606
rect 566 1504 572 1556
rect 624 1544 630 1556
rect 753 1547 811 1553
rect 753 1544 765 1547
rect 624 1516 765 1544
rect 624 1504 630 1516
rect 753 1513 765 1516
rect 799 1513 811 1547
rect 753 1507 811 1513
rect 566 1204 572 1216
rect 527 1176 572 1204
rect 566 1164 572 1176
rect 624 1164 630 1216
rect 201 1114 2382 1136
rect 201 1062 234 1114
rect 286 1062 298 1114
rect 350 1062 1234 1114
rect 1286 1062 1298 1114
rect 1350 1062 2234 1114
rect 2286 1062 2298 1114
rect 2350 1062 2382 1114
rect 201 1040 2382 1062
rect 887 887 2289 893
rect 887 853 899 887
rect 933 876 1067 887
rect 933 853 940 876
rect 887 847 940 853
rect 566 796 572 808
rect 527 768 572 796
rect 566 756 572 768
rect 624 756 630 808
rect 934 715 940 847
rect 887 709 940 715
rect 887 675 899 709
rect 933 684 940 709
rect 992 853 1067 876
rect 1101 853 1235 887
rect 1269 853 1403 887
rect 1437 853 1571 887
rect 1605 853 1739 887
rect 1773 853 1907 887
rect 1941 853 2075 887
rect 2109 853 2243 887
rect 2277 853 2289 887
rect 992 847 2289 853
rect 992 715 998 847
rect 992 709 2289 715
rect 992 684 1067 709
rect 933 675 1067 684
rect 1101 675 1235 709
rect 1269 675 1403 709
rect 1437 675 1571 709
rect 1605 675 1739 709
rect 1773 675 1907 709
rect 1941 675 2075 709
rect 2109 675 2243 709
rect 2277 675 2289 709
rect 887 669 2289 675
rect 201 570 2382 592
rect 201 518 734 570
rect 786 518 798 570
rect 850 518 1734 570
rect 1786 518 1798 570
rect 1850 518 2382 570
rect 201 496 2382 518
<< via1 >>
rect 234 2150 286 2202
rect 298 2150 350 2202
rect 1234 2150 1286 2202
rect 1298 2150 1350 2202
rect 2234 2150 2286 2202
rect 2298 2150 2350 2202
rect 572 1887 624 1896
rect 572 1853 581 1887
rect 581 1853 615 1887
rect 615 1853 624 1887
rect 572 1844 624 1853
rect 1400 1797 1452 1940
rect 1400 1768 1403 1797
rect 1403 1768 1437 1797
rect 1437 1768 1452 1797
rect 734 1606 786 1658
rect 798 1606 850 1658
rect 1734 1606 1786 1658
rect 1798 1606 1850 1658
rect 572 1504 624 1556
rect 572 1207 624 1216
rect 572 1173 581 1207
rect 581 1173 615 1207
rect 615 1173 624 1207
rect 572 1164 624 1173
rect 234 1062 286 1114
rect 298 1062 350 1114
rect 1234 1062 1286 1114
rect 1298 1062 1350 1114
rect 2234 1062 2286 1114
rect 2298 1062 2350 1114
rect 572 799 624 808
rect 572 765 581 799
rect 581 765 615 799
rect 615 765 624 799
rect 572 756 624 765
rect 940 684 992 876
rect 734 518 786 570
rect 798 518 850 570
rect 1734 518 1786 570
rect 1798 518 1850 570
<< metal2 >>
rect 224 2204 360 2213
rect 280 2202 304 2204
rect 286 2150 298 2202
rect 280 2148 304 2150
rect 224 2139 360 2148
rect 1224 2204 1360 2213
rect 1280 2202 1304 2204
rect 1286 2150 1298 2202
rect 1280 2148 1304 2150
rect 1224 2139 1360 2148
rect 2224 2204 2360 2213
rect 2280 2202 2304 2204
rect 2286 2150 2298 2202
rect 2280 2148 2304 2150
rect 2224 2139 2360 2148
rect 1400 1940 1452 1946
rect 572 1896 624 1902
rect 572 1838 624 1844
rect 584 1562 612 1838
rect 1400 1762 1452 1768
rect 724 1660 860 1669
rect 780 1658 804 1660
rect 786 1606 798 1658
rect 780 1604 804 1606
rect 724 1595 860 1604
rect 572 1556 624 1562
rect 572 1498 624 1504
rect 1008 1480 1064 1489
rect 1412 1487 1440 1762
rect 1724 1660 1860 1669
rect 1780 1658 1804 1660
rect 1786 1606 1798 1658
rect 1780 1604 1804 1606
rect 1724 1595 1860 1604
rect 1412 1460 1564 1487
rect 1412 1459 1508 1460
rect 1008 1255 1064 1264
rect 1508 1255 1564 1264
rect 952 1227 1064 1255
rect 572 1216 624 1222
rect 572 1158 624 1164
rect 224 1116 360 1125
rect 280 1114 304 1116
rect 286 1062 298 1114
rect 280 1060 304 1062
rect 224 1051 360 1060
rect 584 814 612 1158
rect 952 882 980 1227
rect 1224 1116 1360 1125
rect 1280 1114 1304 1116
rect 1286 1062 1298 1114
rect 1280 1060 1304 1062
rect 1224 1051 1360 1060
rect 2224 1116 2360 1125
rect 2280 1114 2304 1116
rect 2286 1062 2298 1114
rect 2280 1060 2304 1062
rect 2224 1051 2360 1060
rect 940 876 992 882
rect 572 808 624 814
rect 572 750 624 756
rect 940 678 992 684
rect 724 572 860 581
rect 780 570 804 572
rect 786 518 798 570
rect 780 516 804 518
rect 724 507 860 516
rect 1724 572 1860 581
rect 1780 570 1804 572
rect 1786 518 1798 570
rect 1780 516 1804 518
rect 1724 507 1860 516
<< via2 >>
rect 224 2202 280 2204
rect 304 2202 360 2204
rect 224 2150 234 2202
rect 234 2150 280 2202
rect 304 2150 350 2202
rect 350 2150 360 2202
rect 224 2148 280 2150
rect 304 2148 360 2150
rect 1224 2202 1280 2204
rect 1304 2202 1360 2204
rect 1224 2150 1234 2202
rect 1234 2150 1280 2202
rect 1304 2150 1350 2202
rect 1350 2150 1360 2202
rect 1224 2148 1280 2150
rect 1304 2148 1360 2150
rect 2224 2202 2280 2204
rect 2304 2202 2360 2204
rect 2224 2150 2234 2202
rect 2234 2150 2280 2202
rect 2304 2150 2350 2202
rect 2350 2150 2360 2202
rect 2224 2148 2280 2150
rect 2304 2148 2360 2150
rect 724 1658 780 1660
rect 804 1658 860 1660
rect 724 1606 734 1658
rect 734 1606 780 1658
rect 804 1606 850 1658
rect 850 1606 860 1658
rect 724 1604 780 1606
rect 804 1604 860 1606
rect 1008 1264 1064 1480
rect 1724 1658 1780 1660
rect 1804 1658 1860 1660
rect 1724 1606 1734 1658
rect 1734 1606 1780 1658
rect 1804 1606 1850 1658
rect 1850 1606 1860 1658
rect 1724 1604 1780 1606
rect 1804 1604 1860 1606
rect 1508 1264 1564 1460
rect 224 1114 280 1116
rect 304 1114 360 1116
rect 224 1062 234 1114
rect 234 1062 280 1114
rect 304 1062 350 1114
rect 350 1062 360 1114
rect 224 1060 280 1062
rect 304 1060 360 1062
rect 1224 1114 1280 1116
rect 1304 1114 1360 1116
rect 1224 1062 1234 1114
rect 1234 1062 1280 1114
rect 1304 1062 1350 1114
rect 1350 1062 1360 1114
rect 1224 1060 1280 1062
rect 1304 1060 1360 1062
rect 2224 1114 2280 1116
rect 2304 1114 2360 1116
rect 2224 1062 2234 1114
rect 2234 1062 2280 1114
rect 2304 1062 2350 1114
rect 2350 1062 2360 1114
rect 2224 1060 2280 1062
rect 2304 1060 2360 1062
rect 724 570 780 572
rect 804 570 860 572
rect 724 518 734 570
rect 734 518 780 570
rect 804 518 850 570
rect 850 518 860 570
rect 724 516 780 518
rect 804 516 860 518
rect 1724 570 1780 572
rect 1804 570 1860 572
rect 1724 518 1734 570
rect 1734 518 1780 570
rect 1804 518 1850 570
rect 1850 518 1860 570
rect 1724 516 1780 518
rect 1804 516 1860 518
<< metal3 >>
rect 202 2204 382 2224
rect 202 2148 224 2204
rect 280 2148 304 2204
rect 360 2148 382 2204
rect 202 1116 382 2148
rect 202 1060 224 1116
rect 280 1060 304 1116
rect 360 1060 382 1116
rect 202 496 382 1060
rect 702 1660 882 2224
rect 702 1604 724 1660
rect 780 1604 804 1660
rect 860 1604 882 1660
rect 702 572 882 1604
rect 982 1480 1102 2224
rect 982 1264 1008 1480
rect 1064 1264 1102 1480
rect 982 1239 1102 1264
rect 1202 2204 1382 2224
rect 1202 2148 1224 2204
rect 1280 2148 1304 2204
rect 1360 2148 1382 2204
rect 702 516 724 572
rect 780 516 804 572
rect 860 516 882 572
rect 702 496 882 516
rect 1202 1116 1382 2148
rect 1482 1460 1602 2224
rect 1482 1264 1508 1460
rect 1564 1264 1602 1460
rect 1482 1239 1602 1264
rect 1702 1660 1882 2224
rect 1702 1604 1724 1660
rect 1780 1604 1804 1660
rect 1860 1604 1882 1660
rect 1202 1060 1224 1116
rect 1280 1060 1304 1116
rect 1360 1060 1382 1116
rect 1202 496 1382 1060
rect 1702 572 1882 1604
rect 1702 516 1724 572
rect 1780 516 1804 572
rect 1860 516 1882 572
rect 1702 496 1882 516
rect 2202 2204 2382 2224
rect 2202 2148 2224 2204
rect 2280 2148 2304 2204
rect 2360 2148 2382 2204
rect 2202 1116 2382 2148
rect 2202 1060 2224 1116
rect 2280 1060 2304 1116
rect 2360 1060 2382 1116
rect 2202 496 2382 1060
use sky130_fd_sc_hd__buf_16  const_one_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701272208
transform 1 0 276 0 1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701272208
transform -1 0 828 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_16  const_zero_buf
timestamp 1701272208
transform 1 0 276 0 1 544
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701272208
transform -1 0 1196 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1701272208
transform -1 0 552 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  sky130_fd_sc_hd__decap_12_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701272208
transform -1 0 2392 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701272208
transform 1 0 2300 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1701272208
transform 1 0 2300 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1701272208
transform 1 0 184 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_0
timestamp 1701272208
transform 1 0 1196 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1
timestamp 1701272208
transform 1 0 184 0 1 1632
box -38 -48 130 592
<< labels >>
flabel metal3 s 1202 496 1382 2224 0 FreeSans 960 90 0 0 vccd
port 1 nsew power bidirectional
flabel metal3 s 2202 496 2382 2224 0 FreeSans 960 90 0 0 vccd
port 1 nsew power bidirectional
flabel metal3 s 1702 496 1882 2224 0 FreeSans 960 90 0 0 vssd
port 2 nsew ground bidirectional
flabel metal3 s 702 496 882 2224 0 FreeSans 960 90 0 0 vssd
port 2 nsew ground bidirectional
flabel metal3 s 202 496 382 2224 0 FreeSans 960 90 0 0 vccd
port 1 nsew power bidirectional
flabel metal3 s 982 1424 1102 2224 0 FreeSans 480 90 0 0 zero
port 3 nsew signal tristate
flabel metal3 s 1482 1424 1602 2224 0 FreeSans 480 90 0 0 one
port 0 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 2800 2600
<< end >>
