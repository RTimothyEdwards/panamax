magic
tech sky130A
magscale 1 2
timestamp 1725852642
<< checkpaint >>
rect -1260 27307 2636 42471
rect -1260 13482 2635 27307
rect -1260 13468 2636 13482
rect -1260 13433 2996 13468
rect -1268 13425 2996 13433
rect -1447 13126 2996 13425
rect -1821 12852 2996 13126
rect -1821 12677 3019 12852
rect -2158 10305 3019 12677
rect -2158 9143 2998 10305
rect -2158 1871 2996 9143
rect -2158 -1041 3852 1871
rect -2158 -1274 2996 -1041
rect -2158 -1676 2674 -1274
rect -2158 -1827 2075 -1676
rect -2158 -2276 1738 -1827
<< metal2 >>
rect 496 1100 624 1114
rect 496 609 511 1100
rect 610 609 624 1100
rect 496 0 624 609
rect 752 1100 880 1114
rect 752 609 767 1100
rect 866 609 880 1100
rect 752 0 880 609
<< via2 >>
rect 511 609 610 1100
rect 767 609 866 1100
<< metal3 >>
rect 496 12221 624 12222
rect 0 12177 624 12221
rect 0 11684 71 12177
rect 564 11684 624 12177
rect 0 11627 624 11684
rect 15 11538 302 11565
rect 15 11367 58 11538
rect 266 11367 302 11538
rect 15 11330 302 11367
rect 15 611 156 11330
rect 496 1100 624 11627
rect 496 609 511 1100
rect 610 609 624 1100
rect 496 594 624 609
rect 752 11268 880 12222
rect 1423 11548 1738 11565
rect 1423 11354 1453 11548
rect 1714 11354 1738 11548
rect 1423 11329 1738 11354
rect 752 11220 1375 11268
rect 752 10727 813 11220
rect 1306 10727 1375 11220
rect 752 10674 1375 10727
rect 752 1100 880 10674
rect 1589 10552 1738 11329
rect 752 609 767 1100
rect 866 609 880 1100
rect 1212 10403 1738 10552
rect 1212 611 1361 10403
rect 752 594 880 609
<< via3 >>
rect 71 11684 564 12177
rect 58 11367 266 11538
rect 1453 11354 1714 11548
rect 813 10727 1306 11220
<< metal4 >>
rect 0 12177 624 12221
rect 0 11684 71 12177
rect 564 11684 624 12177
rect 0 11627 624 11684
rect 15 11538 302 11565
rect 15 11367 58 11538
rect 266 11367 302 11538
rect 15 11330 302 11367
rect 1423 11548 1738 11565
rect 1423 11354 1453 11548
rect 1714 11354 1738 11548
rect 1423 11329 1738 11354
rect 752 11220 1376 11268
rect 752 10727 813 11220
rect 1306 10727 1376 11220
rect 752 10674 1376 10727
<< labels >>
flabel metal2 s 752 0 880 609 0 FreeSans 960 270 0 0 amuxbus_b_n
port 0 nsew
flabel metal2 s 496 0 624 609 0 FreeSans 960 270 0 0 amuxbus_a_n
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 1375 41000
string flatten true
<< end >>
