* NGSPICE file created from panamax.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_16 A VGND VNB VPB VPWR X
X0 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X35 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X36 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X39 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X40 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X41 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X42 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X43 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
X0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
.ends

.subckt constant_block one vccd zero vssd
Xconst_zero_buf const_source/LO vssd vssd vccd vccd zero sky130_fd_sc_hd__buf_16
Xconst_source vssd vssd vccd vccd const_source/HI const_source/LO sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_12_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xconst_one_buf const_source/HI vssd vssd vccd vccd one sky130_fd_sc_hd__buf_16
Xsky130_fd_sc_hd__decap_4_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
.ends

.subckt chip_io_ovt_connects_horiz one zero m2_266_24343# m2_548_2675# m2_744_19814#
+ m2_640_5575# constant_block_0/vccd VSUBS
Xconstant_block_0 one constant_block_0/vccd zero VSUBS constant_block
.ends

* Black-box entry subcircuit for sky130_fd_io__top_gpio_ovtv2 abstract view
.subckt sky130_fd_io__top_gpio_ovtv2 VSSIO_Q VSWITCH VSSIO VSSD VSSA VDDIO_Q VDDIO
+ VDDA VCCHIB VCCD PAD AMUXBUS_A AMUXBUS_B DM[0] DM[1] DM[2] INP_DIS VTRIP_SEL IB_MODE_SEL[0]
+ IB_MODE_SEL[1] SLEW_CTL[0] SLEW_CTL[1] HYS_TRIM HLD_OVR ENABLE_H HLD_H_N ENABLE_VDDA_H
+ ANALOG_EN ENABLE_INP_H IN IN_H VINREF OUT ANALOG_POL ANALOG_SEL SLOW OE_N TIE_HI_ESD
+ TIE_LO_ESD PAD_A_ESD_0_H PAD_A_ESD_1_H PAD_A_NOESD_H ENABLE_VSWITCH_H ENABLE_VDDIO
.ends

.subckt sky130_fd_io__com_ctl_ls_octl VCC_IO VPB OUT_H_N OUT_H IN RST_H SET_H HLD_H_N
+ a_992_934# a_181_1305# a_n17_1379#
X0 a_361_1391# a_181_1305# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# a_181_1305# a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_634_829# a_992_934# a_181_1305# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X7 a_361_1391# a_181_1305# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X8 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X17 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=1
X18 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_181_1305# IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X20 a_957_1391# a_181_1305# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X22 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X23 a_n17_1379# IN a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X24 a_724_1391# a_181_1305# a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X26 a_957_1391# a_181_1305# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X27 a_634_829# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X28 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X29 a_724_1391# a_181_1305# a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_128_1391# a_181_1305# a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X31 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_octl DM_H[1] DM_H[0] DM_H[2] DM_H_N[0] DM_H_N[1] DM_H_N[2]
+ PUEN_2OR1_H PDEN_H_N[1] PDEN_H_N[0] SLOW SLOW_H VCC_IO a_n8755_2384# a_n9051_2020#
+ w_n9346_2317# a_n9227_2020# a_n9283_2046# a_5840_3586# m1_n8913_3102# VPWR a_n8875_2020#
+ a_4338_3622# a_3924_6676# a_n8931_2384# a_4514_3388# SLOW_H_N VGND a_5813_4576#
+ HLD_I_H_N OD_H
Xsky130_fd_io__com_ctl_ls_octl_0 VCC_IO VPWR SLOW_H_N SLOW_H SLOW OD_H VGND HLD_I_H_N
+ m2_5755_2254# VPWR VGND sky130_fd_io__com_ctl_ls_octl
X0 a_n8755_2384# a_n9280_2384# a_n8755_2046# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X1 a_n9107_2384# a_n9227_2020# a_n9280_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X2 VCC_IO DM_H_N[0] a_4520_6066# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X3 a_3871_7368# a_3924_6676# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X4 a_4634_3414# a_4514_3388# a_4458_3414# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X5 a_4872_6702# DM_H_N[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X6 VCC_IO DM_H[2] a_3966_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X7 a_4996_5728# a_4520_6066# PUEN_2OR1_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X8 VCC_IO a_4347_7368# a_5651_5728# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X9 a_5813_4576# a_5693_4550# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X10 VCC_IO a_5052_5702# PUEN_2OR1_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X11 a_5488_3924# DM_H_N[1] a_5315_3924# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X12 VCC_IO a_5720_3560# a_5840_3586# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X13 VCC_IO DM_H[0] a_5052_5702# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X14 a_4282_3816# DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X15 VCC_IO DM_H_N[0] a_5175_7368# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X16 a_4634_3816# a_3933_3414# a_4458_3414# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X17 a_4491_4619# a_4371_4587# a_4315_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X18 PDEN_H_N[1] a_5651_6702# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X19 a_5315_3924# DM_H_N[1] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X20 a_5513_4576# a_3871_7368# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X21 VCC_IO DM_H[1] a_4667_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X22 a_4044_6066# DM_H_N[1] a_3871_6066# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X23 a_n8931_2384# a_n9051_2020# a_n9107_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X24 a_n8755_2046# a_n8875_2020# a_n9283_2046# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X25 PDEN_H_N[0] a_5651_5728# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X26 a_4520_6066# a_3871_6066# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X27 a_4347_7368# DM_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X28 a_n8931_2384# a_n9280_2384# a_n8755_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X29 VCC_IO a_4458_3414# a_5488_3924# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X30 a_5513_4576# a_3871_7368# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.1855 ps=1.93 w=0.7 l=0.6
X31 a_4371_4587# DM_H[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X32 VGND a_4458_3414# a_5315_3924# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X33 VCC_IO a_5693_4550# a_5813_4576# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X34 a_4338_3622# DM_H[0] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X35 PUEN_2OR1_H a_4520_6066# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X36 VGND PUEN_2OR1_H a_4044_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X37 PDEN_H_N[1] a_5651_6702# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X38 a_5348_7368# a_4872_6702# a_5175_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X39 VCC_IO DM_H_N[0] a_4520_6066# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X40 VGND a_5651_6702# PDEN_H_N[1] VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X41 VCC_IO DM_H[1] a_4347_7368# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X42 a_5840_3586# a_5720_3560# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X43 VCC_IO DM_H_N[1] a_4872_6702# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X44 a_n8755_2384# a_n8875_2020# a_n8931_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X45 VCC_IO a_4347_7368# a_5651_5728# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X46 a_4458_3414# a_4338_3622# a_4282_3816# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X47 a_4338_3622# DM_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X48 a_4315_5349# DM_H[2] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X49 VCC_IO a_5175_7368# a_5651_6702# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X50 a_4667_5349# a_4371_4587# a_4491_4619# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X51 VGND DM_H_N[2] a_3871_6066# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X52 VGND a_5693_4550# a_5813_4576# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X53 a_5840_3586# a_5720_3560# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X54 a_5813_4576# a_5693_4550# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X55 a_5348_5728# a_4491_4619# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X56 VGND a_5651_5728# PDEN_H_N[0] VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X57 VGND a_3933_3414# a_4634_3414# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X58 a_4315_4619# DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X59 a_5693_4550# a_5513_4576# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X60 a_4667_4619# a_3966_4619# a_4491_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X61 PDEN_H_N[0] a_5651_5728# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X62 a_4044_6066# DM_H_N[1] a_3871_6066# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X63 VGND DM_H_N[0] a_5348_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X64 a_3871_7368# a_3924_6676# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X65 a_4872_6702# DM_H_N[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X66 VCC_IO a_5720_3560# a_5840_3586# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X67 a_4282_3816# DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X68 VCC_IO DM_H[0] a_4634_3816# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X69 VCC_IO PUEN_2OR1_H a_3871_7368# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X70 a_4634_3816# a_3933_3414# a_4458_3414# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X71 a_5813_4576# a_5693_4550# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X72 a_4491_4619# DM_H[1] a_4315_5349# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X73 a_n9280_2384# a_n9227_2020# a_n9283_2046# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X74 VGND a_3966_4619# a_4667_5349# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X75 a_5175_7368# a_4872_6702# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X76 VGND a_5720_3560# a_5840_3586# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X77 VGND a_5052_5702# a_4996_5728# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X78 VCC_IO a_5651_6702# PDEN_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X79 a_5052_5702# DM_H[0] a_5348_5728# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X80 a_n8931_2384# a_n9280_2384# a_n8755_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X81 VGND DM_H[2] a_3933_3414# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X82 a_5720_3560# a_5315_3924# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X83 a_4491_4619# a_4371_4587# a_4315_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X84 VCC_IO DM_H[1] a_4667_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X85 a_4520_7368# DM_H[0] a_4347_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X86 VCC_IO DM_H[2] a_3966_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X87 PUEN_2OR1_H a_4520_6066# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X88 VCC_IO DM_H[2] a_3933_3414# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X89 VCC_IO DM_H_N[2] a_4044_6066# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X90 a_n9283_2046# a_n9051_2020# a_n9280_2384# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X91 a_4371_4587# DM_H[1] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X92 a_5052_5702# a_4491_4619# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X93 a_4520_5728# a_3871_6066# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X94 VCC_IO DM_H_N[0] a_5175_7368# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X95 VCC_IO a_5651_5728# PDEN_H_N[0] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X96 a_n8755_2384# a_n8875_2020# a_n8931_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X97 a_5488_3924# DM_H_N[1] a_5315_3924# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X98 a_4371_4587# DM_H[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X99 VGND DM_H[1] a_4520_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X100 a_n9107_2384# a_n9227_2020# a_n9280_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X101 a_4872_6702# DM_H_N[1] a_4872_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X102 VGND a_5175_7368# a_5651_6702# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X103 a_5693_4550# a_5513_4576# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X104 PDEN_H_N[0] a_5651_5728# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X105 PDEN_H_N[1] a_5651_6702# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X106 a_4338_3622# DM_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X107 VCC_IO a_5052_5702# PUEN_2OR1_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X108 a_4347_7368# DM_H[0] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X109 a_4520_6066# DM_H_N[0] a_4520_5728# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X110 VCC_IO DM_H[0] a_5052_5702# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X111 a_5513_4576# a_3871_7368# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X112 VGND a_4347_7368# a_5651_5728# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X113 a_n8931_2384# a_n9051_2020# a_n9107_2384# w_n9346_2317# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X114 VCC_IO a_4458_3414# a_5488_3924# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X115 a_4044_7368# a_3924_6676# a_3871_7368# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X116 a_4872_7368# DM_H_N[2] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X117 a_5693_4550# a_5513_4576# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X118 a_4458_3414# DM_H[0] a_4282_3414# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X119 VCC_IO DM_H[0] a_4634_3816# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X120 VCC_IO DM_H[1] a_4347_7368# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X121 a_4520_6066# a_3871_6066# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X122 a_3871_6066# DM_H_N[1] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X123 VCC_IO DM_H_N[1] a_4872_6702# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X124 VCC_IO a_5175_7368# a_5651_6702# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X125 VCC_IO DM_H_N[2] a_4044_6066# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X126 VCC_IO PUEN_2OR1_H a_3871_7368# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X127 a_5720_3560# a_5315_3924# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X128 VCC_IO a_5693_4550# a_5813_4576# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X129 a_5052_5702# a_4491_4619# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X130 a_5840_3586# a_5720_3560# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X131 a_5175_7368# a_4872_6702# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X132 VCC_IO a_5651_5728# PDEN_H_N[0] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X133 a_4458_3414# a_4338_3622# a_4282_3816# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X134 VCC_IO a_5651_6702# PDEN_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X135 a_4315_4619# DM_H[2] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X136 VGND DM_H[2] a_3966_4619# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X137 a_4667_4619# a_3966_4619# a_4491_4619# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X138 a_5720_3560# a_5315_3924# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X139 a_4282_3414# DM_H[2] VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X140 VCC_IO DM_H[2] a_3933_3414# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
.ends

.subckt sky130_fd_io__gpio_dat_ls_1v2 IN OUT_H_N RST_H SET_H HLD_H_N VCC_IO VGND OUT_H
+ VPWR_KA
X0 a_2251_36# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X1 a_28_633# SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X2 a_1720_1202# HLD_H_N a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.5
X3 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X4 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X5 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X6 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR_KA a_2251_2228# a_2251_36# VPWR_KA sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X11 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X12 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X13 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X14 a_28_633# a_28_14# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X15 VGND IN a_2251_2228# VGND sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X16 OUT_H a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X17 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X18 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X19 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X20 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X21 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X22 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X23 VGND a_28_633# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X24 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X25 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X26 a_2251_2228# IN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X27 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X28 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X29 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X30 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X31 VGND a_28_633# a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X32 a_2251_2228# IN VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X33 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X34 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X35 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X36 a_28_633# a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X37 a_28_14# a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X38 VGND a_2251_2228# a_2251_36# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X39 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X40 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X41 a_1251_128# HLD_H_N a_28_633# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.56 as=1.325 ps=10.53 w=5 l=0.5
X42 VCC_IO a_28_14# OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X43 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X44 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X45 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X46 VGND RST_H a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X47 OUT_H_N a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X48 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X49 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_io__gpio_dat_lsv2 IN OUT_H_N RST_H SET_H HLD_H_N VCC_IO VGND OUT_H
+ VPWR_KA a_28_14#
X0 a_2251_36# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X1 a_28_633# SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X2 a_1720_1202# HLD_H_N a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.5
X3 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X4 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X5 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X6 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR_KA a_2251_2228# a_2251_36# VPWR_KA sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X11 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X12 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X13 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X14 a_28_633# a_28_14# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X15 VGND IN a_2251_2228# VGND sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X16 OUT_H a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X17 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X18 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X19 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X20 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X21 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X22 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X23 VGND a_28_633# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X24 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X25 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X26 a_2251_2228# IN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X27 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X28 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X29 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X30 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X31 VGND a_28_633# a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X32 a_2251_2228# IN VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X33 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X34 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X35 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X36 a_28_633# a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X37 a_28_14# a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X38 VGND a_2251_2228# a_2251_36# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X39 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X40 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X41 a_1251_128# HLD_H_N a_28_633# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.56 as=1.325 ps=10.53 w=5 l=0.5
X42 VCC_IO a_28_14# OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X43 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X44 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X45 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X46 VGND RST_H a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X47 OUT_H_N a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X48 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X49 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_io__com_cclat PU_DIS_H PD_DIS_H VGND OE_H_N DRVHI_H VCC_IO DRVLO_H_N
X0 a_947_1193# DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X1 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X2 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X3 a_3417_1193# DRVHI_H a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X4 a_4762_1193# DRVHI_H a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X5 VGND DRVHI_H a_2361_1095# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X6 VCC_IO PU_DIS_H a_638_279# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X7 VCC_IO a_2361_1095# DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X8 DRVLO_H_N a_2361_1095# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X9 DRVHI_H a_947_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X10 a_2361_1095# DRVHI_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X11 VCC_IO a_947_1193# DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X12 DRVLO_H_N a_2361_1095# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X13 VCC_IO a_2361_1095# DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X14 DRVHI_H a_947_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X15 VCC_IO a_947_1193# DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X16 VGND PU_DIS_H a_638_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X17 a_4762_1193# DRVHI_H a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X18 a_2361_1095# PD_DIS_H a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X19 VGND PD_DIS_H a_2361_1095# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X20 a_505_1193# a_176_279# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X21 a_3417_1193# DRVHI_H a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X22 a_2361_1095# PD_DIS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X23 VCC_IO a_638_279# a_947_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X24 VGND a_947_1193# DRVHI_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X25 DRVLO_H_N a_2361_1095# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X26 VGND a_947_1193# DRVHI_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X27 a_987_279# a_176_279# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X28 DRVHI_H a_947_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X29 a_4762_1193# PD_DIS_H a_2361_1095# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X30 DRVHI_H a_947_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X31 VCC_IO OE_H_N a_176_279# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X32 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X33 a_2361_1095# PD_DIS_H a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X34 a_987_279# DRVLO_H_N a_1628_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X35 VGND a_2361_1095# DRVLO_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X36 a_947_1193# a_176_279# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X37 DRVHI_H a_947_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X38 VGND OE_H_N a_176_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X39 VCC_IO a_947_1193# DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X40 VCC_IO a_2361_1095# DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X41 DRVLO_H_N a_2361_1095# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X42 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X43 DRVHI_H a_947_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X44 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.6
X45 a_4762_1193# PD_DIS_H a_2361_1095# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X46 VGND a_947_1193# DRVHI_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X47 VGND a_176_279# a_987_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X48 a_947_1193# a_638_279# a_1628_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X49 VGND a_2361_1095# DRVLO_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X50 DRVLO_H_N a_2361_1095# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X51 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X52 a_505_1193# a_176_279# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X53 a_1628_279# DRVLO_H_N a_987_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X54 DRVLO_H_N a_2361_1095# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X55 VGND a_505_1193# a_2361_1095# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X56 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X57 VGND a_176_279# a_987_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X58 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X59 VGND a_2361_1095# DRVLO_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X60 a_2361_1095# a_505_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X61 a_987_279# a_176_279# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X62 a_1628_279# a_638_279# a_947_1193# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
.ends

.subckt sky130_fd_io__com_opath_datoev2 OE_H DRVLO_H_N VCC_IO HLD_I_OVR_H a_5565_99#
+ OUT OE_N sky130_fd_io__com_cclat_0/PD_DIS_H VPWR_KA DRVHI_H li_5565_99# sky130_fd_io__gpio_dat_ls_1v2_0/SET_H
+ VGND OD_H
Xsky130_fd_io__gpio_dat_ls_1v2_0 OUT sky130_fd_io__com_cclat_0/PU_DIS_H VGND sky130_fd_io__gpio_dat_ls_1v2_0/SET_H
+ HLD_I_OVR_H VCC_IO VGND sky130_fd_io__com_cclat_0/PD_DIS_H VPWR_KA sky130_fd_io__gpio_dat_ls_1v2
Xsky130_fd_io__gpio_dat_lsv2_0 OE_N OE_H VGND OD_H HLD_I_OVR_H VCC_IO VGND sky130_fd_io__com_cclat_0/OE_H_N
+ VPWR_KA a_28_1762# sky130_fd_io__gpio_dat_lsv2
Xsky130_fd_io__com_cclat_0 sky130_fd_io__com_cclat_0/PU_DIS_H sky130_fd_io__com_cclat_0/PD_DIS_H
+ VGND sky130_fd_io__com_cclat_0/OE_H_N DRVHI_H VCC_IO DRVLO_H_N sky130_fd_io__com_cclat
.ends

.subckt sky130_fd_io__com_pdpredrvr_weakv2 DRVLO_H_N PDEN_H_N VGND_IO VCC_IO PD_H
X0 PD_H DRVLO_H_N a_73_866# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X1 a_73_866# PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X2 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X3 VGND_IO DRVLO_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X4 VCC_IO PDEN_H_N a_73_866# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_octl_mux SEL_H_N A_H Y_H B_H SEL_H a_1266_1185# w_1191_2415#
X0 Y_H SEL_H A_H a_1266_1185# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X1 A_H SEL_H_N Y_H w_1191_2415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X2 Y_H SEL_H B_H w_1191_2415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X3 B_H SEL_H_N Y_H a_1266_1185# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_pdpredrvr_strong sky130_fd_io__gpiov2_octl_mux_0/SEL_H
+ sky130_fd_io__gpiov2_octl_mux_0/B_H sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N sky130_fd_io__gpiov2_octl_mux_0/w_1191_2415#
+ sky130_fd_io__gpiov2_octl_mux_0/A_H sky130_fd_io__gpiov2_octl_mux_0/Y_H VSUBS
Xsky130_fd_io__gpiov2_octl_mux_0 sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N sky130_fd_io__gpiov2_octl_mux_0/A_H
+ sky130_fd_io__gpiov2_octl_mux_0/Y_H sky130_fd_io__gpiov2_octl_mux_0/B_H sky130_fd_io__gpiov2_octl_mux_0/SEL_H
+ VSUBS sky130_fd_io__gpiov2_octl_mux_0/w_1191_2415# sky130_fd_io__gpiov2_octl_mux
.ends

.subckt sky130_fd_io__feascom_pupredrvr_nbiasv2 EN_H EN_H_N VGND_IO DRVHI_H NBIAS
+ PUEN_H VCC_IO PU_H_N a_261_220# a_2821_220# a_2874_118# a_1772_220#
X0 VCC_IO a_250_1898# a_1507_1397# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X1 VGND_IO a_261_220# a_261_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X2 a_1507_1397# a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X3 a_261_220# a_261_220# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X4 a_1672_194# a_207_1014# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X5 NBIAS a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.1925 ps=1.385 w=1 l=0.8
X6 a_250_1898# a_562_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X7 VGND_IO a_1672_194# a_1772_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X8 VCC_IO a_250_1898# a_2874_118# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X9 NBIAS NBIAS a_261_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X10 VGND_IO a_1672_194# a_1772_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R0 a_562_1898# m1_2838_1831# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R1 m1_1014_127# NBIAS sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X11 VCC_IO DRVHI_H a_562_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.185 pd=1.515 as=0.14 ps=1.28 w=1 l=0.5
R2 m1_1014_800# NBIAS sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X12 a_261_220# a_261_220# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R3 m1_575_1252# EN_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X13 a_250_1898# DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X14 VGND_IO DRVHI_H a_207_1014# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.32375 pd=2.015 as=0.265 ps=2.53 w=1 l=0.6
X15 VGND_IO a_207_1014# NBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R4 m1_2838_1794# a_620_1263# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R5 m1_612_1252# a_620_1263# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X16 VGND_IO a_250_1898# a_1004_990# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=4
X17 NBIAS NBIAS a_261_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X18 VCC_IO a_250_1898# NBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X19 a_2874_118# a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.0375 ps=5.515 w=5 l=0.5
X20 a_583_914# EN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.2025 pd=1.77 as=0.32375 ps=2.015 w=1.5 l=0.5
X21 a_2821_220# a_2874_118# a_2874_118# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X22 a_1772_220# a_1672_194# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R6 m1_1409_1332# NBIAS sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X23 NBIAS a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
R7 m1_1608_646# a_1772_220# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X24 a_207_1014# DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X25 a_250_1898# a_562_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X26 a_261_220# NBIAS NBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X27 NBIAS EN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X28 VCC_IO a_250_1898# a_1507_1397# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.8
X29 a_2821_220# a_2821_220# a_1672_194# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X30 VCC_IO a_562_1898# a_250_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.0375 pd=5.515 as=0.42 ps=3.28 w=3 l=0.5
X31 a_1772_220# a_1672_194# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R8 m1_2596_1928# a_2421_2014# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X32 a_1507_1397# a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
R9 m1_2596_1928# a_250_1898# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X33 VCC_IO EN_H a_250_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X34 a_562_1898# PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X35 a_2421_2014# PU_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.185 ps=1.515 w=0.42 l=8
R10 m1_702_1715# PU_H_N sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R11 m1_1409_1332# a_1507_1397# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X36 VCC_IO a_250_1898# NBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X37 a_737_914# a_620_1263# a_583_914# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.2025 pd=1.77 as=0.2025 ps=1.77 w=1.5 l=0.5
X38 a_261_220# NBIAS NBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X39 VGND_IO a_261_220# a_261_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R12 m1_1014_800# a_1004_990# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R13 m1_1046_126# a_261_220# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X40 VCC_IO a_562_1898# a_250_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R14 a_620_1263# m1_702_1715# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X41 a_250_1898# DRVHI_H a_737_914# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.2025 ps=1.77 w=1.5 l=0.5
R15 m1_1608_646# a_261_220# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X42 a_1672_194# a_2821_220# a_2821_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X43 a_562_1898# a_620_1263# a_620_1263# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X44 a_1672_194# VCC_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=8
X45 VCC_IO DRVHI_H a_207_1014# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1925 pd=1.385 as=0.14 ps=1.28 w=1 l=0.5
X46 a_2874_118# a_2874_118# a_2821_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_pupredrvr_strong_nd2 DRVHI_H PUEN_H EN_FAST[0] EN_FAST[1]
+ EN_FAST[2] EN_FAST[3] VGND_IO VCC_IO PU_H_N a_158_632#
X0 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.6
X1 a_311_632# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.1575 pd=1.71 as=0.3975 ps=3.53 w=1.5 l=0.5
X2 VGND_IO EN_FAST[3] a_311_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.1575 ps=1.71 w=1.5 l=1
R0 PU_H_N m1_1184_866# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X3 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X4 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.6
R1 m1_1184_866# a_158_632# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X5 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X6 a_158_632# DRVHI_H a_809_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.165 ps=1.72 w=1.5 l=0.5
X7 a_1008_2434# PU_H_N sky130_fd_pr__res_generic_po w=0.33 l=4
X8 a_809_632# EN_FAST[2] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.165 pd=1.72 as=0.21 ps=1.78 w=1.5 l=1
X9 a_158_632# DRVHI_H a_809_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.165 ps=1.72 w=1.5 l=0.5
X10 a_1008_2434# a_158_632# sky130_fd_pr__res_generic_po w=0.33 l=11
X11 a_311_1060# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.1575 pd=1.71 as=0.3975 ps=3.53 w=1.5 l=0.5
X12 VGND_IO EN_FAST[0] a_311_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.1575 ps=1.71 w=1.5 l=1
X13 PU_H_N DRVHI_H a_158_109# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
X14 VGND_IO PUEN_H a_158_109# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
X15 a_809_1060# EN_FAST[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.165 pd=1.72 as=0.21 ps=1.78 w=1.5 l=1
.ends

.subckt sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a DRVHI_H PUEN_H EN_FAST[0] EN_FAST[1]
+ EN_FAST[2] EN_FAST[3] VGND_IO VCC_IO PU_H_N a_353_606# a_609_606#
X0 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.6
X1 a_311_632# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.1575 pd=1.71 as=0.3975 ps=3.53 w=1.5 l=0.5
X2 VGND_IO a_353_606# a_311_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.1575 ps=1.71 w=1.5 l=1
R0 PU_H_N m1_1184_866# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X3 VGND_IO PUEN_H a_158_199# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
X4 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X5 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.6
R1 m1_1184_866# a_158_632# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X6 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X7 a_158_632# DRVHI_H a_809_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.165 ps=1.72 w=1.5 l=0.5
X8 a_1008_2434# PU_H_N sky130_fd_pr__res_generic_po w=0.33 l=4
X9 a_809_632# a_609_606# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.165 pd=1.72 as=0.21 ps=1.78 w=1.5 l=1
X10 a_158_632# DRVHI_H a_809_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.165 ps=1.72 w=1.5 l=0.5
X11 a_1008_2434# a_158_632# sky130_fd_pr__res_generic_po w=0.33 l=11
X12 a_311_1060# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.1575 pd=1.71 as=0.3975 ps=3.53 w=1.5 l=0.5
X13 VGND_IO EN_FAST[0] a_311_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.1575 ps=1.71 w=1.5 l=1
X14 PU_H_N DRVHI_H a_158_199# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
X15 a_809_1060# EN_FAST[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.165 pd=1.72 as=0.21 ps=1.78 w=1.5 l=1
.ends

.subckt sky130_fd_io__gpio_pupredrvr_strongv2 VCC_IO PU_H_N[3] PUEN_H PU_H_N[2] SLOW_H_N
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220# DRVHI_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ VSUBS
Xsky130_fd_io__feascom_pupredrvr_nbiasv2_0 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VSUBS DRVHI_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ PUEN_H VCC_IO PU_H_N[2] sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2
Xsky130_fd_io__gpiov2_pupredrvr_strong_nd2_0 DRVHI_H PUEN_H sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[0]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[1] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[2]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] VSUBS VCC_IO PU_H_N[3] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2
Xsky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0 DRVHI_H PUEN_H sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] VSUBS VCC_IO PU_H_N[2]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a
R0 m1_4655_1468# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X0 VCC_IO PUEN_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
R1 m1_6555_1273# VSUBS sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R2 m1_6556_1365# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[0] sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X1 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N SLOW_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
R3 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[1] m1_6299_1273# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R4 VSUBS m1_6266_605# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R5 m1_5759_509# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R6 m1_4777_1326# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R7 m1_5786_421# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R8 m1_4655_1468# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R9 m1_6266_568# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[2] sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R10 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] m1_5786_421# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X2 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
R11 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] m1_6300_1402# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R12 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[2] m1_6265_477# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R13 m1_5722_509# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R14 m1_6300_1365# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[1] sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R15 m1_6299_1273# VSUBS sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R16 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[0] m1_6555_1273# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R17 m1_6265_477# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X3 VSUBS PUEN_H a_483_1179# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X4 a_483_1179# SLOW_H_N sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X5 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VSUBS VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
R18 m1_4740_1326# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R19 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] m1_6556_1402# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
.ends

.subckt sky130_fd_io__gpiov2_obpredrvr sky130_fd_io__gpio_pupredrvr_strongv2_0/SLOW_H_N
+ sky130_fd_io__com_pdpredrvr_weakv2_0/PDEN_H_N sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N
+ sky130_fd_io__com_pdpredrvr_weakv2_0/VCC_IO sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/A_H sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H sky130_fd_io__com_pdpredrvr_weakv2_0/PD_H
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/DRVHI_H sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/PU_H_N[2] sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/w_1191_2415#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/PU_H_N[3] sky130_fd_io__com_pdpredrvr_weakv2_0/DRVLO_H_N
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/B_H sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ VSUBS sky130_fd_io__gpio_pupredrvr_strongv2_0/VCC_IO
Xsky130_fd_io__com_pdpredrvr_weakv2_0 sky130_fd_io__com_pdpredrvr_weakv2_0/DRVLO_H_N
+ sky130_fd_io__com_pdpredrvr_weakv2_0/PDEN_H_N VSUBS sky130_fd_io__com_pdpredrvr_weakv2_0/VCC_IO
+ sky130_fd_io__com_pdpredrvr_weakv2_0/PD_H sky130_fd_io__com_pdpredrvr_weakv2
Xsky130_fd_io__gpiov2_pdpredrvr_strong_0 sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/B_H sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/w_1191_2415#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/A_H sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ VSUBS sky130_fd_io__gpiov2_pdpredrvr_strong
Xsky130_fd_io__gpio_pupredrvr_strongv2_0 sky130_fd_io__gpio_pupredrvr_strongv2_0/VCC_IO
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/PU_H_N[3] sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/PU_H_N[2] sky130_fd_io__gpio_pupredrvr_strongv2_0/SLOW_H_N
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/DRVHI_H sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ VSUBS sky130_fd_io__gpio_pupredrvr_strongv2
.ends

.subckt sky130_fd_io__gpiov2_octl_dat VPWR_KA VGND SLOW HLD_I_OVR_H OD_H SLOW_H_N
+ DRVHI_H PU_H_N[2] PU_H_N[1] PU_H_N[0] PD_H[1] PD_H[0] PD_H[4] PD_H[3] PD_H[2] a_1106_3203#
+ a_3125_3203# a_4416_3253# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ a_n433_1745# a_8354_4056# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ DM_H[0] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ DM_H[1] DM_H_N[0] DM_H_N[1] DM_H[2] DM_H_N[2] a_1415_3203# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ OE_N sky130_fd_io__com_opath_datoev2_0/li_5565_99# a_9656_1708# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ HLD_I_H_N a_1528_3203# a_2205_3177# VGND_IO VPWR sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ OUT VCC_IO PU_H_N[3]
Xsky130_fd_io__gpiov2_octl_0 DM_H[1] DM_H[0] DM_H[2] DM_H_N[0] DM_H_N[1] DM_H_N[2]
+ sky130_fd_io__gpiov2_octl_0/PUEN_2OR1_H sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1]
+ sky130_fd_io__gpiov2_octl_0/PDEN_H_N[0] SLOW sky130_fd_io__gpiov2_octl_0/SLOW_H
+ VCC_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N
+ DM_H[1] VCC_IO DM_H[0] VGND a_7799_1681# VCC_IO VPWR DM_H[2] a_13335_4479# VCC_IO
+ VCC_IO a_13335_4479# SLOW_H_N VGND sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H
+ HLD_I_H_N OD_H sky130_fd_io__gpiov2_octl
Xsky130_fd_io__com_opath_datoev2_0 sky130_fd_io__com_opath_datoev2_0/OE_H DRVLO_H_N
+ VCC_IO HLD_I_OVR_H VGND OUT OE_N sky130_fd_io__com_opath_datoev2_0/sky130_fd_io__com_cclat_0/PD_DIS_H
+ VPWR_KA DRVHI_H sky130_fd_io__com_opath_datoev2_0/li_5565_99# OD_H VGND OD_H sky130_fd_io__com_opath_datoev2
Xsky130_fd_io__gpiov2_obpredrvr_0 SLOW_H_N sky130_fd_io__gpiov2_octl_0/PDEN_H_N[0]
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N
+ VCC_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/A_H
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H
+ PD_H[0] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ DRVHI_H sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ PU_H_N[2] VCC_IO PU_H_N[3] DRVLO_H_N DRVLO_H_N sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ VGND_IO VCC_IO sky130_fd_io__gpiov2_obpredrvr
X0 a_8354_4056# PD_H[4] a_8354_3203# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
X1 a_3125_3203# a_1415_3203# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R0 a_7638_3476# m1_8994_2579# sky130_fd_pr__res_generic_m1 w=2.5 l=10m
X2 a_1528_3203# a_2205_3177# a_2205_3177# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X3 a_1415_3203# a_1528_3203# a_1528_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X4 VCC_IO a_1415_3203# a_3125_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X5 VCC_IO DRVLO_H_N a_1159_3105# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X6 VGND_IO a_7610_2597# a_1106_3203# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=1
X7 PU_H_N[0] a_7799_1681# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.6
X8 a_2205_3177# a_2205_3177# a_1528_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R1 a_10919_675# m1_10778_2585# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X9 a_1528_3203# a_1528_3203# a_1415_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X10 VGND_IO a_7799_1681# a_7743_1707# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X11 VCC_IO a_4416_3253# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X12 a_11758_843# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=2
X13 sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X14 VCC_IO DRVHI_H PU_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X15 PD_H[3] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X16 a_1106_3203# a_1106_3203# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X17 a_4416_3253# a_4416_3253# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X18 VCC_IO a_n461_1863# a_9290_3718# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X19 VGND PD_H[4] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/A_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.5
X20 a_1415_3203# a_1159_3105# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
R2 m1_10510_2769# a_7462_4229# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X21 a_7161_3177# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.335 ps=2.67 w=1 l=0.6
X22 PD_H[3] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H a_11053_559# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.5
X23 VCC_IO DRVHI_H PU_H_N[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X24 a_n408_4001# sky130_fd_io__gpiov2_octl_0/SLOW_H a_n112_4027# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X25 VCC_IO a_7610_2597# a_8026_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
X26 a_7462_4229# a_7161_3177# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.21 ps=1.42 w=1 l=0.6
X27 a_9290_3718# a_1106_3203# a_9882_3718# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
R3 m1_8330_3159# a_7610_2597# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R4 m1_10378_2704# m1_10351_2626# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X28 a_10564_1155# a_11085_1123# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X29 a_n408_1837# sky130_fd_io__gpiov2_octl_0/SLOW_H a_n112_1863# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X30 a_8876_944# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X31 VCC_IO sky130_fd_io__gpiov2_octl_0/SLOW_H a_n408_1837# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
R5 m1_10312_2627# a_1106_3203# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R6 m1_8994_2542# a_7512_2477# sky130_fd_pr__res_generic_m1 w=2.5 l=10m
R7 m1_7727_3684# a_7462_4229# sky130_fd_pr__res_generic_m1 w=0.64 l=10m
X32 VCC_IO a_n461_4027# a_9935_2938# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.63 pd=3.42 as=0.42 ps=3.28 w=3 l=0.6
R8 a_8354_3203# m1_8330_3159# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R9 m1_10312_2627# m1_10351_2626# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R10 a_7462_4229# m1_10378_2741# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X33 a_4416_3253# a_1106_3203# a_1106_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X34 a_7512_2477# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X35 a_11053_559# a_10919_675# a_10398_443# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.5
X36 a_1106_3203# a_1106_3203# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R11 m1_10523_1531# VCC_IO sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X37 a_1106_3203# a_1106_3203# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X38 a_9656_1708# DRVHI_H PU_H_N[1] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X39 a_3125_3203# a_1415_3203# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X40 a_4416_3253# a_1106_3203# a_1106_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X41 PD_H[2] DRVLO_H_N a_10194_3718# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X42 a_12137_3347# DRVLO_H_N PD_H[4] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=1
R12 m1_9138_2849# a_1106_3203# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X43 a_1159_3105# DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X44 VGND a_n408_4001# a_n461_4027# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X45 PD_H[3] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X46 VCC_IO sky130_fd_io__gpiov2_octl_0/SLOW_H a_n408_4001# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X47 VGND_IO a_7610_2597# a_9179_2770# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=1
X48 PD_H[3] sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X49 VCC_IO a_1415_3203# a_3125_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X50 a_3125_3203# a_1415_3203# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X51 a_7613_3603# a_7462_4229# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.315 pd=3.21 as=0.795 ps=6.53 w=3 l=0.5
R13 a_11085_1123# m1_10523_1531# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X52 sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X53 VCC_IO a_1159_3105# a_1106_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X54 a_10873_1155# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X55 PD_H[2] DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X56 VGND a_n408_1837# a_n461_1863# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X57 VCC_IO a_n408_1837# a_n461_1863# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X58 a_11862_3305# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_11009_3305# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
X59 PD_H[3] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H a_10564_1155# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X60 a_8876_944# DRVLO_H_N PD_H[1] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X61 PD_H[4] sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X62 a_7755_3603# a_7638_3476# a_7613_3603# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.315 pd=3.21 as=0.315 ps=3.21 w=3 l=0.5
X63 PD_H[2] DRVLO_H_N a_9882_3718# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X64 VCC_IO PD_H[4] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/A_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
R14 m1_10547_2769# a_10919_675# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X65 sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.1855 ps=1.93 w=0.7 l=0.6
X66 a_11009_3305# DRVLO_H_N PD_H[2] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
X67 a_9656_1708# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X68 a_n112_4027# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X69 VGND_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X70 VCC_IO sky130_fd_io__gpiov2_octl_0/SLOW_H a_n408_1837# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X71 a_7610_2597# DRVLO_H_N a_7755_3603# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.315 ps=3.21 w=3 l=0.5
X72 VGND_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
R15 m1_4181_3684# a_4416_3253# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X73 a_n112_1863# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X74 a_9179_2770# a_7610_2597# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=1
X75 VGND_IO DRVLO_H_N PD_H[2] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X76 VGND_IO a_n461_4027# a_7161_3177# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.42 as=0.14 ps=1.28 w=1 l=0.6
X77 a_n408_1837# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X78 VGND_IO sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] PD_H[2] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X79 VCC_IO a_n408_4001# a_n461_4027# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X80 a_4416_3253# a_4416_3253# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X81 a_1106_3203# a_7610_2597# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=1
X82 a_8354_4056# PD_H[4] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
R16 m1_7764_3684# a_7638_3476# sky130_fd_pr__res_generic_m1 w=0.64 l=10m
X83 a_4416_3253# a_1106_3203# a_1106_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X84 a_1528_3203# a_2205_3177# a_2205_3177# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X85 a_1106_3203# a_1106_3203# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X86 a_10194_3718# DRVLO_H_N PD_H[2] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R17 m1_5837_4210# a_1106_3203# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X87 PU_H_N[1] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X88 a_1415_3203# a_1528_3203# a_1528_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X89 a_7638_3476# a_7638_3476# a_7512_2477# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X90 a_2205_3177# a_2205_3177# a_1528_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X91 VGND_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/PUEN_H a_9656_1708# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X92 a_1106_3203# a_7161_3177# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X93 PU_H_N[0] DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.6
X94 VGND_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X95 VCC_IO a_4416_3253# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X96 VCC_IO a_4416_3253# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R18 m1_9138_2849# a_9179_2770# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X97 a_4416_3253# a_4416_3253# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X98 a_9290_3718# a_n461_1863# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X99 VCC_IO sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_11009_3747# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
X100 PU_H_N[1] DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X101 VCC_IO a_n408_1837# a_n461_1863# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X102 VCC_IO sky130_fd_io__gpiov2_octl_0/SLOW_H a_n408_4001# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X103 a_n408_4001# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X104 VGND_IO DRVLO_H_N a_7512_2477# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X105 VCC_IO a_1106_3203# a_12137_3347# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=1
R19 m1_10375_2471# a_1106_3203# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R20 m1_4181_3684# a_3125_3203# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X106 PD_H[3] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H a_10849_843# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=2
X107 VCC_IO VGND_IO a_1415_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=8
R21 m1_8014_3310# a_8026_3203# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X108 VGND_IO sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] PD_H[3] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X109 a_7610_2597# a_7512_2477# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.6
X110 a_10398_443# a_n461_1863# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X111 a_4416_3253# a_1106_3203# a_1106_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R22 m1_10375_2471# a_10919_675# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R23 m1_9297_3844# PD_H[4] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X112 a_10398_443# a_11085_1123# a_11053_559# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.5
X113 a_n408_1837# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X114 VGND_IO DRVLO_H_N a_1159_3105# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X115 VGND_IO DRVLO_H_N PD_H[4] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X116 PD_H[2] a_n461_1863# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X117 VCC_IO DRVHI_H PU_H_N[0] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X118 PD_H[1] sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X119 VGND_IO DRVLO_H_N a_7610_2597# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X120 a_11862_3305# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_9290_3718# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
X121 VCC_IO a_1415_3203# a_3125_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X122 a_4416_3253# a_4416_3253# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
R24 a_1106_3203# m1_8014_3310# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X123 VCC_IO a_1415_3203# a_3125_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X124 a_9290_3718# a_n461_1863# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X125 a_3125_3203# a_1415_3203# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X126 a_9935_2938# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_7161_3177# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=1.005 ps=6.67 w=3 l=0.6
X127 VCC_IO a_n408_4001# a_n461_4027# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X128 a_1528_3203# a_1528_3203# a_1415_3203# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R25 m1_9297_3844# a_7638_3476# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X129 a_11053_559# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.5
X130 VCC_IO a_10919_675# a_10873_1155# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X131 a_7462_4229# a_7161_3177# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.63 ps=3.42 w=3 l=0.6
R26 m1_5874_4210# a_4416_3253# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X132 a_10398_443# sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_11758_843# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=2
X133 VCC_IO a_4416_3253# a_4416_3253# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X134 a_10194_3718# a_1106_3203# a_9290_3718# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X135 PU_H_N[1] DRVHI_H a_9656_1708# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X136 PD_H[1] DRVLO_H_N a_8876_944# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X137 a_7610_2597# a_7462_4229# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X138 VGND_IO DRVLO_H_N PD_H[1] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X139 a_7743_1707# DRVHI_H PU_H_N[0] VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X140 PD_H[4] DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X141 a_2205_3177# a_7610_2597# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.6
R27 m1_10778_2548# a_11085_1123# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X142 a_9882_3718# DRVLO_H_N PD_H[2] VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X143 VCC_IO sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_10849_843# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
X144 PD_H[4] DRVLO_H_N a_11009_3747# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=4
X145 a_n408_4001# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/SEL_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X146 PD_H[4] DRVLO_H_N a_12137_3347# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X147 VCC_IO a_n461_1863# a_10398_443# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X148 VCC_IO sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] a_8876_944# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
.ends

.subckt sky130_fd_io__com_res_weak_bentbigres a_419_6804# a_419_8054# a_n256_8772#
+ a_419_8146# a_n258_6046# a_419_9396# a_n2_6046#
X0 a_419_8054# a_419_6804# sky130_fd_pr__res_generic_po w=0.8 l=6
X1 a_n256_8772# a_n258_6046# sky130_fd_pr__res_generic_po w=0.8 l=12
X2 a_419_9396# a_419_8146# sky130_fd_pr__res_generic_po w=0.8 l=6
X3 a_n258_6046# a_n2_6046# sky130_fd_pr__res_generic_po w=0.8 l=50
.ends

.subckt sky130_fd_io__com_res_weak RA RB sky130_fd_io__com_res_weak_bentbigres_0/a_n258_6046#
+ a_n160_10423# li_n135_8054# li_n135_6820# a_n160_9488#
Xsky130_fd_io__com_res_weak_bentbigres_0 li_n135_6820# li_n135_8054# li_n135_6820#
+ li_n135_8054# sky130_fd_io__com_res_weak_bentbigres_0/a_n258_6046# a_n160_9488#
+ RA sky130_fd_io__com_res_weak_bentbigres
R0 m1_n147_9555# a_n160_9488# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R1 m1_n146_7434# li_n135_6820# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
X0 a_n160_10423# a_n160_9838# sky130_fd_pr__res_generic_po w=0.8 l=1.5
X1 a_n160_9838# a_n160_9488# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R2 a_n160_10423# m1_n147_10115# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R3 a_n160_9488# m1_n147_8777# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R4 a_n160_10423# m1_532_10115# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R5 a_517_9818# m1_532_9534# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R6 m1_n147_8777# li_n135_8054# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R7 m1_n147_10115# a_n160_9838# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R8 m1_532_10115# a_517_9818# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
X2 a_517_9818# RB sky130_fd_pr__res_generic_po w=0.8 l=1.5
R9 m1_532_9534# RB sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R10 a_n160_9838# m1_n147_9555# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R11 li_n135_8054# m1_n146_7735# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
X3 a_n160_10423# a_517_9818# sky130_fd_pr__res_generic_po w=0.8 l=1.5
.ends

.subckt sky130_fd_io__pfet_con_diff_wo_abt_270v2 w_415_600# a_2303_1380# a_13777_1380#
+ a_8817_1380# a_4287_1380# a_7263_1380# a_12223_1380# a_9247_1380# a_2865_1380# a_5841_1380#
+ a_4849_1380# a_10801_1380# a_14135_1380# a_1311_1380# a_12785_1380# a_7825_1380#
+ a_3295_1380# a_9809_1380# a_1001_1552# a_6271_1380# a_5279_1380# a_11231_1380# a_10239_1380#
+ a_8255_1380# a_1873_1380# a_13215_1380# a_3857_1380# a_11793_1380# a_881_1380# a_6833_1380#
X0 a_1001_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.975 pd=6.19 as=3.775 ps=11.51 w=5 l=0.6
X1 w_415_600# a_10239_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X2 a_1001_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X3 a_1001_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X4 w_415_600# a_14135_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.72 as=2.975 ps=6.19 w=5 l=0.6
X5 w_415_600# a_3295_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X6 a_1001_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X7 w_415_600# a_2303_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X8 w_415_600# a_7263_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X9 a_1001_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X10 w_415_600# a_11231_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X11 a_1001_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X12 w_415_600# a_10239_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X13 a_1001_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X14 w_415_600# a_3295_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X15 w_415_600# a_2303_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X16 w_415_600# a_7263_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X17 a_1001_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X18 a_1001_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X19 a_1001_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X20 w_415_600# a_13215_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X21 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X22 w_415_600# a_6271_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X23 a_1001_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X24 w_415_600# a_5279_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X25 a_1001_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X26 a_1001_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X27 a_1001_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X28 w_415_600# a_13215_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X29 w_415_600# a_9247_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X30 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X31 w_415_600# a_6271_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X32 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=4.325 ps=11.73 w=5 l=0.6
X33 w_415_600# a_5279_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X34 a_1001_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X35 a_1001_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X36 a_1001_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X37 w_415_600# a_9247_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X38 a_1001_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X39 w_415_600# a_12223_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X40 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=4.325 ps=11.73 w=5 l=0.6
X41 a_1001_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X42 a_1001_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X43 w_415_600# a_4287_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X44 a_1001_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X45 w_415_600# a_8255_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X46 w_415_600# a_12223_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X47 a_1001_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.975 pd=6.19 as=3.775 ps=11.51 w=5 l=0.6
X48 a_1001_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X49 a_1001_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X50 w_415_600# a_4287_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X51 w_415_600# a_14135_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.72 as=2.975 ps=6.19 w=5 l=0.6
X52 a_1001_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X53 w_415_600# a_11231_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X54 w_415_600# a_8255_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X55 a_1001_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpio_pudrvr_strongv2 PU_H_N[3] PU_H_N[2] VCC_IO m1_1330_n459#
+ TIE_HI_ESD m1_6027_281# m1_3418_50# VNB a_14575_n157# m1_6652_281# m1_3028_333#
+ PAD m1_14880_n614# li_9083_n155#
Xsky130_fd_io__pfet_con_diff_wo_abt_270v2_0 VCC_IO PU_H_N[2] m1_14229_1478# m1_8837_1478#
+ PU_H_N[3] PU_H_N[3] m1_11745_1478# m1_8837_1478# PU_H_N[2] PU_H_N[3] PU_H_N[3] m1_10391_1478#
+ m1_14229_1478# PU_H_N[2] PU_H_N[2] PU_H_N[3] PU_H_N[2] m1_10391_1478# PAD PU_H_N[3]
+ PU_H_N[3] m1_11745_1478# m1_10391_1478# m1_8837_1478# PU_H_N[2] m1_13667_1478# PU_H_N[3]
+ m1_11745_1478# PU_H_N[2] PU_H_N[3] sky130_fd_io__pfet_con_diff_wo_abt_270v2
R0 m2_14075_657# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R1 m1_14229_1478# m2_14532_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 m1_13667_1478# m2_13593_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R3 m2_12849_n185# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 m1_8837_1478# m2_10673_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 m1_10391_1478# m2_10945_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R6 m2_10673_n208# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 m2_11422_n209# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 m1_13667_1478# m2_14075_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 m2_10197_n209# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 m2_10945_n209# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 m1_11745_1478# m2_12608_116# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 m1_10391_1478# m2_11422_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 m1_11745_1478# m2_12849_116# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 m2_12608_n185# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 m2_13837_658# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 m2_14769_657# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 m2_11186_n208# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R18 m2_14286_658# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X0 TIE_HI_ESD a_14575_n157# sky130_fd_pr__res_generic_po w=0.5 l=10.2
R19 m1_8837_1478# m2_10197_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m1_8837_1478# m2_10439_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 m2_14532_657# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 m1_10391_1478# m2_11186_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R23 m2_13593_657# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 m1_13667_1478# m2_13837_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 m1_14229_1478# m2_14769_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 m1_11745_1478# m2_12365_n184# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 m2_10439_n209# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 m2_12365_n184# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R29 m1_14229_1478# m2_14286_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__nfet_con_diff_wo_abt_270v2 VCC_IO VSSIO PAD a_10282_1285# a_5322_1285#
+ a_12266_1285# a_7306_1285# a_3900_1285# a_2908_1285# a_5884_1285# a_14178_1285#
+ a_10844_1285# a_1354_1285# a_7868_1285# a_12828_1285# a_8860_1285# a_13820_1285#
+ a_4330_1285# a_3338_1285# a_11274_1285# a_6314_1285# a_8298_1285# a_13258_1285#
+ a_9290_1285# a_1916_1285# a_4892_1285# a_6876_1285# a_924_1285# a_11836_1285# a_2346_1285#
+ a_9852_1285#
X0 PAD a_10844_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X1 PAD a_9852_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X2 VSSIO a_2346_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X3 PAD a_1916_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X4 PAD a_6876_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X5 VSSIO a_12266_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X6 VSSIO a_6314_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X7 PAD a_11836_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X8 VSSIO a_9290_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X9 PAD a_4892_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X10 VSSIO a_4330_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X11 PAD a_8860_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X12 VSSIO a_10282_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X13 VSSIO a_3338_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X14 VSSIO a_8298_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X15 PAD a_924_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.425 ps=11.37 w=5 l=0.6
X16 PAD a_3900_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X17 PAD a_13820_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=2.975 pd=6.19 as=3.775 ps=11.51 w=5 l=0.6
X18 PAD a_2908_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X19 PAD a_7868_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X20 VSSIO a_13258_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X21 VSSIO a_7306_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X22 PAD a_12828_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X23 VSSIO a_14178_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.425 pd=11.37 as=2.975 ps=6.19 w=5 l=0.6
X24 VSSIO a_1354_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X25 PAD a_5884_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X26 VSSIO a_11274_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X27 VSSIO a_5322_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X28 PAD a_9852_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X29 PAD a_10844_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X30 VSSIO a_2346_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X31 PAD a_6876_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X32 VSSIO a_6314_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X33 PAD a_1916_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X34 VSSIO a_12266_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X35 PAD a_11836_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X36 PAD a_4892_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X37 VSSIO a_9290_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X38 PAD a_8860_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X39 VSSIO a_10282_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X40 VSSIO a_4330_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X41 PAD a_924_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.425 ps=11.37 w=5 l=0.6
X42 PAD a_3900_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X43 VSSIO a_3338_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X44 VSSIO a_8298_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X45 PAD a_2908_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X46 PAD a_7868_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X47 VSSIO a_7306_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X48 PAD a_13820_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=2.975 pd=6.19 as=3.775 ps=11.51 w=5 l=0.6
X49 VSSIO a_13258_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X50 PAD a_12828_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X51 VSSIO a_1354_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X52 VSSIO a_14178_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.425 pd=11.37 as=2.975 ps=6.19 w=5 l=0.6
X53 PAD a_5884_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X54 VSSIO a_5322_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X55 VSSIO a_11274_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_pddrvr_strong sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_3338_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_4330_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_10282_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_6314_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_12266_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_8298_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_9290_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_1916_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/VSSIO
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_4892_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/VCC_IO
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_10844_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/PAD
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_6876_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_14178_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_2346_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_12828_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_13820_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_924_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_9852_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_5322_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_11274_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_7306_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_13258_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_3900_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_2908_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_5884_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_1354_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_7868_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_11836_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_8860_1285#
Xsky130_fd_io__nfet_con_diff_wo_abt_270v2_0 sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/VCC_IO
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/VSSIO sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/PAD
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_10282_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_5322_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_12266_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_7306_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_3900_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_2908_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_5884_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_14178_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_10844_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_1354_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_7868_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_12828_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_8860_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_13820_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_4330_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_3338_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_11274_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_6314_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_8298_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_13258_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_9290_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_1916_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_4892_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_6876_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_924_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_11836_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_2346_1285# sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/a_9852_1285#
+ sky130_fd_io__nfet_con_diff_wo_abt_270v2
.ends

.subckt sky130_fd_io__com_pudrvr_weakv2 PU_H_N PAD w_258_n30# a_756_297#
X0 PAD PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X1 PAD PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X2 w_258_n30# PU_H_N a_756_297# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X3 w_258_n30# PU_H_N a_756_297# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X4 w_258_n30# PU_H_N PAD w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X5 w_258_n30# PU_H_N PAD w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=1.855 pd=14.53 as=0.98 ps=7.28 w=7 l=0.5
X6 a_756_297# PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X7 a_756_297# PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.855 ps=14.53 w=7 l=0.5
.ends

.subckt sky130_fd_io__res250_sub_small a_10_2# a_2142_2#
X0 a_10_2# a_2142_2# sky130_fd_pr__res_generic_po w=2 l=10.07
.ends

.subckt sky130_fd_io__res250only_small PAD ROUT
Xsky130_fd_io__res250_sub_small_0 PAD ROUT sky130_fd_io__res250_sub_small
.ends

.subckt sky130_fd_io__gpio_pddrvr_weakv2 PD_H PAD dw_n122_84# w_168_168#
X0 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.6
X1 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.6
X2 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.6
X3 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.6
X4 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.6
X5 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpio_odrvr_subv2 VGND PD_H[0] PD_H[2] PD_H[1] PD_H[3] TIE_LO_ESD
+ FORCE_HI_H_N FORCE_LO_H FORCE_LOVOL_H PU_H_N[0] PU_H_N[1] PU_H_N[2] PU_H_N[3] VSSIO_AMX
+ VGND_IO w_588_14893# m3_6107_13425# w_n915_9930# li_5884_n9263# m2_8191_n10933#
+ sky130_fd_io__gpiov2_pddrvr_strong_0/sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/VSSIO
+ sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614# sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ TIE_HI_ESD m1_2782_13727# PAD w_5497_14893# VCC_IO
Xsky130_fd_io__com_res_weak_0 sky130_fd_io__com_res_weak_0/RA sky130_fd_io__com_res_weak_0/RB
+ sky130_fd_io__com_res_weak_0/sky130_fd_io__com_res_weak_bentbigres_0/a_n258_6046#
+ sky130_fd_io__com_res_weak_0/a_n160_10423# sky130_fd_io__com_res_weak_0/li_n135_8054#
+ sky130_fd_io__com_res_weak_0/li_n135_6820# sky130_fd_io__com_res_weak_0/a_n160_9488#
+ sky130_fd_io__com_res_weak
Xsky130_fd_io__gpio_pudrvr_strongv2_0 PU_H_N[3] PU_H_N[2] VCC_IO VCC_IO TIE_HI_ESD
+ VCC_IO PU_H_N[0] VGND VCC_IO VCC_IO VCC_IO PAD sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155# sky130_fd_io__gpio_pudrvr_strongv2
Xsky130_fd_io__gpiov2_pddrvr_strong_0 m1_11278_13727# m1_9854_13727# PD_H[3] m1_8317_13727#
+ m1_2782_13727# PD_H[2] PD_H[3] m1_12832_13727# sky130_fd_io__gpiov2_pddrvr_strong_0/sky130_fd_io__nfet_con_diff_wo_abt_270v2_0/VSSIO
+ m1_9854_13727# VCC_IO PD_H[3] PAD m1_8317_13727# m1_870_13727# m1_12832_13727# m1_2220_13727#
+ m1_870_13727# m1_12832_13727# PD_H[3] m1_9854_13727# PD_H[3] m1_7742_13727# m1_870_13727#
+ m1_11278_13727# m1_11278_13727# m1_8317_13727# m1_12832_13727# PD_H[2] PD_H[3] PD_H[2]
+ sky130_fd_io__gpiov2_pddrvr_strong
Xsky130_fd_io__com_pudrvr_weakv2_0 PU_H_N[0] sky130_fd_io__com_res_weak_0/RA VCC_IO
+ sky130_fd_io__com_res_weak_0/RA sky130_fd_io__com_pudrvr_weakv2
Xsky130_fd_io__res250only_small_0 PAD sky130_fd_io__com_res_weak_0/RB sky130_fd_io__res250only_small
Xsky130_fd_io__gpio_pddrvr_weakv2_0 PD_H[0] sky130_fd_io__com_res_weak_0/RA VCC_IO
+ w_5497_14893# sky130_fd_io__gpio_pddrvr_weakv2
X0 TIE_LO_ESD VGND_IO sky130_fd_pr__res_generic_po w=0.5 l=10.2
R0 PD_H[2] m2_11414_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X1 VCC_IO PU_H_N[1] a_782_15260# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.855 pd=14.53 as=0.98 ps=7.28 w=7 l=0.5
R1 TIE_LO_ESD m2_1933_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 m2_12848_15816# m1_12832_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X2 a_10314_7886# sky130_fd_io__com_res_weak_0/RB sky130_fd_pr__res_generic_po w=2 l=2
R3 m2_982_15816# m1_870_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 PD_H[2] m2_10071_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X3 a_782_15260# PD_H[1] w_588_14893# w_588_14893# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.6
X4 a_782_15260# PU_H_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.855 ps=14.53 w=7 l=0.5
R5 TIE_LO_ESD m2_9451_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X5 a_9612_7886# a_10314_7886# sky130_fd_pr__res_generic_po w=2 l=3
R6 PD_H[3] m2_7318_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 m2_13278_15816# m1_12832_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X6 a_782_15260# PD_H[1] w_588_14893# w_588_14893# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.6
R8 TIE_LO_ESD m2_499_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 PD_H[2] m2_6889_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 m2_11414_15816# m1_11278_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X7 a_782_15260# PD_H[1] w_588_14893# w_588_14893# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.6
R11 m2_1933_15816# m1_2220_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 TIE_LO_ESD m2_10931_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 m2_10071_15816# m1_9854_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 m2_9451_15816# m1_8317_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 PD_H[3] m2_1650_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 m2_7318_15817# m1_7742_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X8 a_782_15260# PU_H_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.855 ps=14.53 w=7 l=0.5
R17 PD_H[2] m2_1345_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R18 m2_499_15816# m1_870_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 m2_6889_15816# m1_7742_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m2_10931_15816# m1_9854_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 TIE_LO_ESD m2_13707_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 m1_9882_7996# a_10314_7886# sky130_fd_pr__res_generic_m1 w=1.32 l=10m
R23 PD_H[3] m2_9020_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 PD_H[3] m2_740_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 m2_1650_15816# m1_2220_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 PD_H[2] m2_8591_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X9 a_782_15260# PU_H_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
R27 m1_9882_7996# a_9612_7886# sky130_fd_pr__res_generic_m1 w=1.32 l=10m
R28 m2_1345_15817# m1_2220_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X10 VCC_IO PU_H_N[1] a_782_15260# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
R29 PD_H[3] m2_10500_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R30 m2_9020_15817# m1_8317_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R31 PD_H[3] m2_11843_15817# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R32 m2_13707_15817# m1_12832_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R33 m2_740_15817# m1_870_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R34 m2_8591_15816# m1_8317_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R35 TIE_LO_ESD m2_12274_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R36 TIE_LO_ESD m2_7749_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X11 a_782_15260# PD_H[1] w_588_14893# w_588_14893# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.6
X12 VCC_IO PU_H_N[1] a_782_15260# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.855 pd=14.53 as=0.98 ps=7.28 w=7 l=0.5
X13 a_782_15260# PU_H_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
R37 m2_10500_15817# m1_9854_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R38 m2_11843_15817# m1_11278_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X14 VCC_IO PU_H_N[1] a_782_15260# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
R39 PD_H[2] m2_982_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R40 PD_H[2] m2_12848_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R41 m2_12274_15816# m1_11278_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R42 m2_7749_15816# m1_7742_13727# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R43 PD_H[3] m2_13278_16117# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X15 a_782_15260# a_9612_7886# sky130_fd_pr__res_generic_po w=2 l=5
.ends

.subckt sky130_fd_io__gpio_odrvrv2 PAD PD_H[0] PD_H[1] PD_H[2] PD_H[3] PU_H_N[0] PU_H_N[1]
+ PU_H_N[2] PU_H_N[3] FORCE_HI_H_N FORCE_LO_H VSSIO_AMX w_n915_9930# FORCE_LOVOL_H
+ sky130_fd_io__gpio_odrvr_subv2_0/m3_6107_13425# TIE_LO_ESD TIE_HI_ESD w_5497_14893#
+ sky130_fd_io__gpio_odrvr_subv2_0/li_5884_n9263# sky130_fd_io__gpio_odrvr_subv2_0/m2_8191_n10933#
+ w_588_14893# sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ sky130_fd_io__gpio_odrvr_subv2_0/m1_2782_13727# VGND VCC_IO VGND_IO
Xsky130_fd_io__gpio_odrvr_subv2_0 VGND PD_H[0] PD_H[2] PD_H[1] PD_H[3] TIE_LO_ESD
+ FORCE_HI_H_N FORCE_LO_H FORCE_LOVOL_H PU_H_N[0] PU_H_N[1] PU_H_N[2] PU_H_N[3] VSSIO_AMX
+ VGND_IO w_588_14893# sky130_fd_io__gpio_odrvr_subv2_0/m3_6107_13425# w_n915_9930#
+ sky130_fd_io__gpio_odrvr_subv2_0/li_5884_n9263# sky130_fd_io__gpio_odrvr_subv2_0/m2_8191_n10933#
+ VGND_IO sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ TIE_HI_ESD sky130_fd_io__gpio_odrvr_subv2_0/m1_2782_13727# PAD w_5497_14893# VCC_IO
+ sky130_fd_io__gpio_odrvr_subv2
.ends

.subckt sky130_fd_io__gpio_opathv2 HLD_I_OVR_H HLD_I_H_N OD_H SLOW VPWR sky130_fd_io__gpiov2_octl_dat_0/a_1528_3203#
+ sky130_fd_io__gpiov2_octl_dat_0/a_2205_3177# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ DM_H[0] DM_H_N[0] sky130_fd_io__gpiov2_octl_dat_0/a_1106_3203# DM_H[2] DM_H_N[1]
+ m1_4747_14860# sky130_fd_io__gpio_odrvrv2_0/sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ TIE_LO_ESD sky130_fd_io__gpiov2_octl_dat_0/a_3125_3203# sky130_fd_io__gpiov2_octl_dat_0/a_4416_3253#
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] m2_2157_n626# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ TIE_HI_ESD m1_5007_14796# DM_H[1] PAD sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpiov2_octl_dat_0/a_8354_4056# DM_H_N[2] sky130_fd_io__gpiov2_octl_dat_0/a_1415_3203#
+ VSSIO_AMX sky130_fd_io__gpiov2_octl_dat_0/a_9656_1708# VPWR_KA OE_N OUT VGND VCC_IO
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ VGND_IO
Xsky130_fd_io__gpiov2_octl_dat_0 VPWR_KA VGND SLOW HLD_I_OVR_H OD_H sky130_fd_io__gpiov2_octl_dat_0/SLOW_H_N
+ sky130_fd_io__gpiov2_octl_dat_0/DRVHI_H sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[1]
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[0] sky130_fd_io__gpio_odrvrv2_0/PD_H[1] sky130_fd_io__gpio_odrvrv2_0/PD_H[0]
+ sky130_fd_io__gpiov2_octl_dat_0/PD_H[4] sky130_fd_io__gpio_odrvrv2_0/PD_H[3] sky130_fd_io__gpio_odrvrv2_0/PD_H[2]
+ sky130_fd_io__gpiov2_octl_dat_0/a_1106_3203# sky130_fd_io__gpiov2_octl_dat_0/a_3125_3203#
+ sky130_fd_io__gpiov2_octl_dat_0/a_4416_3253# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ VGND sky130_fd_io__gpiov2_octl_dat_0/a_8354_4056# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ DM_H[0] sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ DM_H[1] DM_H_N[0] DM_H_N[1] DM_H[2] DM_H_N[2] sky130_fd_io__gpiov2_octl_dat_0/a_1415_3203#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ OE_N VGND sky130_fd_io__gpiov2_octl_dat_0/a_9656_1708# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ HLD_I_H_N sky130_fd_io__gpiov2_octl_dat_0/a_1528_3203# sky130_fd_io__gpiov2_octl_dat_0/a_2205_3177#
+ VGND_IO VPWR sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ OUT VCC_IO sky130_fd_io__gpio_odrvrv2_0/PU_H_N[3] sky130_fd_io__gpiov2_octl_dat
Xsky130_fd_io__gpio_odrvrv2_0 PAD sky130_fd_io__gpio_odrvrv2_0/PD_H[0] sky130_fd_io__gpio_odrvrv2_0/PD_H[1]
+ sky130_fd_io__gpio_odrvrv2_0/PD_H[2] sky130_fd_io__gpio_odrvrv2_0/PD_H[3] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[0]
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[1] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[3]
+ VSSIO_AMX VSSIO_AMX VSSIO_AMX w_n815_25161# VSSIO_AMX VGND_IO TIE_LO_ESD TIE_HI_ESD
+ VGND_IO VGND VGND VGND_IO sky130_fd_io__gpio_odrvrv2_0/sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[1] sky130_fd_io__gpiov2_octl_dat_0/PD_H[4] VGND
+ VCC_IO VGND_IO sky130_fd_io__gpio_odrvrv2
.ends

.subckt sky130_fd_io__amux_switch_1v2b AMUXBUS_HV PG_AMX_VDDA_H_N NG_AMX_VPMP_H NG_PAD_VPMP_H
+ PAD_HV_P0 PAD_HV_P1 PG_PAD_VDDIOQ_H_N PAD_HV_N0 PAD_HV_N1 VDDA VSSD PAD_HV_N2 VDDIO
+ PAD_HV_N3 w_7010_315# w_3919_213#
X0 AMUXBUS_HV NG_AMX_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X1 PAD_HV_N0 NG_PAD_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X2 w_3919_213# PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X3 PAD_HV_N1 NG_PAD_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X4 w_7010_315# NG_PAD_VPMP_H PAD_HV_N2 w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X5 AMUXBUS_HV PG_AMX_VDDA_H_N w_3919_213# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X6 w_3919_213# PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X7 w_3919_213# NG_PAD_VPMP_H PAD_HV_N1 w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.96 pd=14.56 as=1.225 ps=7.35 w=7 l=0.5
X8 PAD_HV_N2 NG_PAD_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X9 w_3919_213# NG_AMX_VPMP_H AMUXBUS_HV w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X10 w_3919_213# PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.225 pd=7.35 as=1.96 ps=14.56 w=7 l=0.5
X11 w_3919_213# NG_PAD_VPMP_H PAD_HV_N0 w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=2.205 ps=14.63 w=7 l=0.5
X12 w_7010_315# NG_AMX_VPMP_H AMUXBUS_HV w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X13 w_7010_315# NG_PAD_VPMP_H PAD_HV_N3 w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X14 w_3919_213# NG_PAD_VPMP_H PAD_HV_N1 w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X15 AMUXBUS_HV NG_AMX_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X16 AMUXBUS_HV NG_AMX_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=2.205 pd=14.63 as=0.98 ps=7.28 w=7 l=0.5
X17 w_3919_213# PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=2.205 ps=14.63 w=7 l=0.5
X18 w_7010_315# NG_AMX_VPMP_H AMUXBUS_HV w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X19 AMUXBUS_HV PG_AMX_VDDA_H_N w_3919_213# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X20 AMUXBUS_HV NG_AMX_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.225 pd=7.35 as=1.96 ps=14.56 w=7 l=0.5
X21 PAD_HV_N3 NG_PAD_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X22 PAD_HV_P1 PG_PAD_VDDIOQ_H_N w_3919_213# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=2.205 pd=14.63 as=0.98 ps=7.28 w=7 l=0.5
X23 PAD_HV_P1 PG_PAD_VDDIOQ_H_N w_3919_213# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X24 PAD_HV_N2 NG_PAD_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=2.205 ps=14.63 w=7 l=0.5
X25 AMUXBUS_HV NG_AMX_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X26 PAD_HV_N3 NG_PAD_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X27 w_3919_213# NG_AMX_VPMP_H AMUXBUS_HV w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X28 PAD_HV_N1 NG_PAD_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X29 w_7010_315# NG_PAD_VPMP_H PAD_HV_N2 w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X30 w_7010_315# NG_AMX_VPMP_H AMUXBUS_HV w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=2.205 pd=14.63 as=0.98 ps=7.28 w=7 l=0.5
X31 w_7010_315# NG_AMX_VPMP_H AMUXBUS_HV w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.225 pd=7.35 as=1.96 ps=14.56 w=7 l=0.5
X32 w_3919_213# PG_PAD_VDDIOQ_H_N PAD_HV_P1 VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X33 w_3919_213# PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.205 pd=14.63 as=0.98 ps=7.28 w=7 l=0.5
X34 PAD_HV_P0 PG_PAD_VDDIOQ_H_N w_3919_213# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.225 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X35 w_3919_213# NG_AMX_VPMP_H AMUXBUS_HV w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X36 w_3919_213# NG_PAD_VPMP_H PAD_HV_N0 w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X37 AMUXBUS_HV NG_AMX_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X38 AMUXBUS_HV NG_AMX_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.225 ps=7.35 w=7 l=0.5
X39 w_7010_315# NG_PAD_VPMP_H PAD_HV_N3 w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=2.205 pd=14.63 as=0.98 ps=7.28 w=7 l=0.5
.ends

.subckt sky130_fd_io__res75only_small PAD ROUT
X0 PAD ROUT sky130_fd_pr__res_generic_po w=2 l=3.15
.ends

.subckt sky130_fd_io__inv_1 VNB VPB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
.ends

.subckt sky130_fd_io__nor2_1 vgnd vpwr A Y B vnb vpb
X0 a_116_368# A vpwr vpb sky130_fd_pr__pfet_01v8_hvt ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X1 Y A vgnd vnb sky130_fd_pr__nfet_01v8 ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2 Y B a_116_368# vpb sky130_fd_pr__pfet_01v8_hvt ad=0.3304 pd=2.83 as=0.1512 ps=1.39 w=1.12 l=0.15
X3 vgnd B Y vnb sky130_fd_pr__nfet_01v8 ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
.ends

.subckt sky130_fd_io__nand2_1 VNB VPB VPWR VGND B Y A
X0 a_117_74# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2 Y A a_117_74# VNB sky130_fd_pr__nfet_01v8 ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
.ends

.subckt sky130_fd_io__gpiov2_amux_decoder sky130_fd_io__inv_1_8/A sky130_fd_io__inv_1_0/Y
+ sky130_fd_io__inv_1_11/A sky130_fd_io__inv_1_2/Y sky130_fd_io__inv_1_13/A sky130_fd_io__nor2_1_0/Y
+ sky130_fd_io__inv_1_4/Y sky130_fd_io__nand2_1_0/Y sky130_fd_io__inv_1_1/A sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__nand2_1_2/Y sky130_fd_io__inv_1_6/Y sky130_fd_io__inv_1_3/A sky130_fd_io__nor2_1_1/B
+ sky130_fd_io__inv_1_8/Y sky130_fd_io__nand2_1_1/B sky130_fd_io__nor2_1_1/A sky130_fd_io__inv_1_11/Y
+ sky130_fd_io__inv_1_5/A sky130_fd_io__nand2_1_1/A sky130_fd_io__nor2_1_3/B sky130_fd_io__nor2_1_3/A
+ sky130_fd_io__inv_1_13/Y sky130_fd_io__nand2_1_3/B sky130_fd_io__inv_1_7/A sky130_fd_io__inv_1_10/A
+ sky130_fd_io__nand2_1_3/A sky130_fd_io__inv_1_1/Y sky130_fd_io__inv_1_12/A sky130_fd_io__inv_1_9/A
+ sky130_fd_io__inv_1_8/VGND sky130_fd_io__inv_1_3/Y sky130_fd_io__inv_1_14/A sky130_fd_io__inv_1_0/A
+ sky130_fd_io__nor2_1_1/Y sky130_fd_io__nand2_1_1/Y sky130_fd_io__inv_1_5/Y sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__nor2_1_3/Y sky130_fd_io__inv_1_2/A sky130_fd_io__nor2_1_0/A sky130_fd_io__inv_1_7/Y
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__nand2_1_3/Y sky130_fd_io__inv_1_10/Y sky130_fd_io__nand2_1_0/B
+ sky130_fd_io__inv_1_4/A sky130_fd_io__nand2_1_0/A sky130_fd_io__nor2_1_2/B sky130_fd_io__inv_1_9/Y
+ sky130_fd_io__nor2_1_2/A sky130_fd_io__inv_1_12/Y sky130_fd_io__inv_1_6/A sky130_fd_io__nand2_1_2/B
+ sky130_fd_io__nand2_1_2/A sky130_fd_io__tap_1_2/VPWR sky130_fd_io__tap_1_1/VGND
+ VSUBS sky130_fd_io__inv_1_14/Y sky130_fd_io__tap_1_2/VPB
Xsky130_fd_io__inv_1_10 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__inv_1_10/Y sky130_fd_io__inv_1_10/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_11 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__inv_1_11/Y sky130_fd_io__inv_1_11/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_12 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__inv_1_8/VGND sky130_fd_io__inv_1_12/Y sky130_fd_io__inv_1_12/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_13 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__inv_1_8/VGND sky130_fd_io__inv_1_13/Y sky130_fd_io__inv_1_13/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_14 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_14/Y sky130_fd_io__inv_1_14/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_0 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_0/Y sky130_fd_io__inv_1_0/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_1 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_1/Y sky130_fd_io__inv_1_1/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_2 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_2/Y sky130_fd_io__inv_1_2/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_3 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_3/Y sky130_fd_io__inv_1_3/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_4 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_4/Y sky130_fd_io__inv_1_4/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_5 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__inv_1_5/Y sky130_fd_io__inv_1_5/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_6 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_1/VGND sky130_fd_io__inv_1_6/Y sky130_fd_io__inv_1_6/A sky130_fd_io__inv_1
Xsky130_fd_io__nor2_1_0 sky130_fd_io__tap_1_1/VGND sky130_fd_io__tap_1_2/VPWR sky130_fd_io__nor2_1_0/A
+ sky130_fd_io__nor2_1_0/Y sky130_fd_io__nor2_1_0/B VSUBS sky130_fd_io__tap_1_2/VPB
+ sky130_fd_io__nor2_1
Xsky130_fd_io__inv_1_7 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__inv_1_7/Y sky130_fd_io__inv_1_7/A sky130_fd_io__inv_1
Xsky130_fd_io__nor2_1_2 sky130_fd_io__tap_1_1/VGND sky130_fd_io__tap_1_2/VPWR sky130_fd_io__nor2_1_2/A
+ sky130_fd_io__nor2_1_2/Y sky130_fd_io__nor2_1_2/B VSUBS sky130_fd_io__tap_1_2/VPB
+ sky130_fd_io__nor2_1
Xsky130_fd_io__nor2_1_1 sky130_fd_io__tap_1_1/VGND sky130_fd_io__tap_1_2/VPWR sky130_fd_io__nor2_1_1/A
+ sky130_fd_io__nor2_1_1/Y sky130_fd_io__nor2_1_1/B VSUBS sky130_fd_io__tap_1_2/VPB
+ sky130_fd_io__nor2_1
Xsky130_fd_io__nor2_1_3 sky130_fd_io__tap_1_1/VGND sky130_fd_io__tap_1_2/VPWR sky130_fd_io__nor2_1_3/A
+ sky130_fd_io__nor2_1_3/Y sky130_fd_io__nor2_1_3/B VSUBS sky130_fd_io__tap_1_2/VPB
+ sky130_fd_io__nor2_1
Xsky130_fd_io__inv_1_8 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__inv_1_8/VGND sky130_fd_io__inv_1_8/Y sky130_fd_io__inv_1_8/A sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_9 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__inv_1_9/Y sky130_fd_io__inv_1_9/A sky130_fd_io__inv_1
Xsky130_fd_io__nand2_1_0 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__nand2_1_0/B sky130_fd_io__nand2_1_0/Y sky130_fd_io__nand2_1_0/A
+ sky130_fd_io__nand2_1
Xsky130_fd_io__nand2_1_1 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__inv_1_8/VGND sky130_fd_io__nand2_1_1/B sky130_fd_io__nand2_1_1/Y sky130_fd_io__nand2_1_1/A
+ sky130_fd_io__nand2_1
Xsky130_fd_io__nand2_1_2 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__nand2_1_2/B sky130_fd_io__nand2_1_2/Y sky130_fd_io__nand2_1_2/A
+ sky130_fd_io__nand2_1
Xsky130_fd_io__nand2_1_3 VSUBS sky130_fd_io__tap_1_2/VPB sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__tap_1_2/VGND sky130_fd_io__nand2_1_3/B sky130_fd_io__nand2_1_3/Y sky130_fd_io__nand2_1_3/A
+ sky130_fd_io__nand2_1
.ends

.subckt sky130_fd_io__gpiov2_amux_ctl_logic sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VPWR
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPB sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VPB sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VGND
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_1/VGND sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/VGND
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A VSUBS sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VGND
Xsky130_fd_io__gpiov2_amux_decoder_0 sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/VGND
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VGND
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/B sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPWR sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_1/VGND
+ VSUBS sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPB
+ sky130_fd_io__gpiov2_amux_decoder
.ends

.subckt sky130_fd_io__gpiov2_amux sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_P0 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__res75only_small_0/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N3 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/A
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N2 sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N1 sky130_fd_io__res75only_small_7/ROUT
+ sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N0 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B
+ sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/A
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_P1 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/A
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_P0 sky130_fd_io__res75only_small_13/PAD
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N sky130_fd_io__res75only_small_2/PAD
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/Y
+ sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ sky130_fd_io__amux_switch_1v2b_1/VDDA sky130_fd_io__res75only_small_8/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A
+ sky130_fd_io__res75only_small_9/PAD sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/Y
+ sky130_fd_io__res75only_small_13/ROUT sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y
+ sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H sky130_fd_io__res75only_small_1/PAD
+ sky130_fd_io__res75only_small_8/PAD sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__res75only_small_10/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VPWR
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/B
+ sky130_fd_io__res75only_small_0/PAD sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/A
+ sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_1/VGND
+ sky130_fd_io__res75only_small_9/ROUT w_8674_6609# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__amux_switch_1v2b_0/AMUXBUS_HV sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VPB
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N3 sky130_fd_io__res75only_small_6/ROUT
+ sky130_fd_io__res75only_small_7/PAD sky130_fd_io__amux_switch_1v2b_1/AMUXBUS_HV
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/B
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N2 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N1 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/A
+ w_11765_6609# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y
+ w_8674_4393# w_11765_4495# sky130_fd_io__res75only_small_3/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VGND
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VGND
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N0 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/A
+ sky130_fd_io__amux_switch_1v2b_0/VDDIO sky130_fd_io__res75only_small_5/PAD sky130_fd_io__amux_switch_1v2b_0/PAD_HV_P1
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPB
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/VGND
+ sky130_fd_io__amux_switch_1v2b_1/VDDIO VSUBS
Xsky130_fd_io__amux_switch_1v2b_0 sky130_fd_io__amux_switch_1v2b_0/AMUXBUS_HV sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N
+ sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_P0 sky130_fd_io__amux_switch_1v2b_0/PAD_HV_P1
+ sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N0
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N1 sky130_fd_io__amux_switch_1v2b_1/VDDA
+ VSUBS sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N2 sky130_fd_io__amux_switch_1v2b_0/VDDIO
+ sky130_fd_io__amux_switch_1v2b_0/PAD_HV_N3 w_11765_6609# w_8674_6609# sky130_fd_io__amux_switch_1v2b
Xsky130_fd_io__amux_switch_1v2b_1 sky130_fd_io__amux_switch_1v2b_1/AMUXBUS_HV sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N
+ sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_P0 sky130_fd_io__amux_switch_1v2b_1/PAD_HV_P1
+ sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N0
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N1 sky130_fd_io__amux_switch_1v2b_1/VDDA
+ VSUBS sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N2 sky130_fd_io__amux_switch_1v2b_1/VDDIO
+ sky130_fd_io__amux_switch_1v2b_1/PAD_HV_N3 w_11765_4495# w_8674_4393# sky130_fd_io__amux_switch_1v2b
Xsky130_fd_io__res75only_small_10 sky130_fd_io__res75only_small_10/PAD sky130_fd_io__res75only_small_10/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_11 sky130_fd_io__res75only_small_2/PAD sky130_fd_io__res75only_small_10/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_13 sky130_fd_io__res75only_small_13/PAD sky130_fd_io__res75only_small_13/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_12 sky130_fd_io__res75only_small_1/PAD sky130_fd_io__res75only_small_13/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_0 sky130_fd_io__res75only_small_0/PAD sky130_fd_io__res75only_small_0/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_1 sky130_fd_io__res75only_small_1/PAD sky130_fd_io__res75only_small_3/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_2 sky130_fd_io__res75only_small_2/PAD sky130_fd_io__res75only_small_0/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_3 sky130_fd_io__res75only_small_3/PAD sky130_fd_io__res75only_small_3/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_4 sky130_fd_io__res75only_small_5/PAD sky130_fd_io__res75only_small_4/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__gpiov2_amux_ctl_logic_0 sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_0/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VPWR
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_10/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_2/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPB
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/B
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VPB
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__tap_1_0/VGND
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_1/VGND
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/VGND
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_3/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VPWR
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ VSUBS sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__tap_1_2/VGND
+ sky130_fd_io__gpiov2_amux_ctl_logic
Xsky130_fd_io__res75only_small_5 sky130_fd_io__res75only_small_5/PAD sky130_fd_io__res75only_small_5/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_6 sky130_fd_io__res75only_small_8/PAD sky130_fd_io__res75only_small_6/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_7 sky130_fd_io__res75only_small_7/PAD sky130_fd_io__res75only_small_7/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_8 sky130_fd_io__res75only_small_8/PAD sky130_fd_io__res75only_small_8/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_9 sky130_fd_io__res75only_small_9/PAD sky130_fd_io__res75only_small_9/ROUT
+ sky130_fd_io__res75only_small
.ends

.subckt sky130_fd_io__gpiov2_ipath_hvls OUT OUT_B MODE_NORMAL_N IN_VCCHIB INB_VCCHIB
+ IN_VDDIO MODE_VCCHIB_N MODE_NORMAL MODE_VCCHIB VDDIO_Q VSSD
X0 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X1 a_1752_1955# a_1175_2172# OUT_B VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X2 a_602_2876# IN_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X3 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X4 a_1930_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X5 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X6 a_621_2778# MODE_VCCHIB_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X7 a_2024_2876# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X8 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X9 VDDIO_Q MODE_VCCHIB_N a_1290_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X10 a_1930_201# IN_VCCHIB a_602_2876# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X11 a_621_2778# INB_VCCHIB a_881_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X12 a_881_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X13 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X14 VSSD MODE_VCCHIB a_1752_1955# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X15 VSSD MODE_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X16 VSSD MODE_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X17 a_621_2778# a_602_2876# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X18 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X19 a_1290_2876# a_1175_2172# OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X20 VDDIO_Q MODE_NORMAL_N a_2024_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X21 a_1752_2267# MODE_NORMAL VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X22 a_881_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X23 a_881_201# INB_VCCHIB a_621_2778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X24 a_1175_2172# a_602_2876# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.3975 ps=3.53 w=1.5 l=0.5
X25 VDDIO_Q MODE_NORMAL a_2911_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X26 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X27 VSSD MODE_VCCHIB a_881_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X28 VDDIO_Q a_621_2778# a_602_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X29 a_2024_2876# IN_VDDIO OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X30 OUT_B a_1175_2172# a_1290_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X31 OUT_B IN_VDDIO a_1752_2267# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X32 VSSD MODE_VCCHIB a_881_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X33 a_881_201# INB_VCCHIB a_621_2778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X34 a_602_2876# IN_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X35 a_2911_2876# MODE_VCCHIB OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X36 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X37 a_1930_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X38 a_1175_2172# a_602_2876# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.3975 ps=3.53 w=1.5 l=0.5
X39 a_1290_2876# MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X40 OUT_B IN_VDDIO a_2024_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_vcchib_in_buf IN_H MODE_VCCHIB_LV_N VCCHIB VSSD OUT OUT_N
X0 VCCHIB MODE_VCCHIB_LV_N a_612_2476# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.25
X1 a_612_2476# MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.25
X2 VCCHIB MODE_VCCHIB_LV_N a_612_2476# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.25
X3 a_538_595# a_591_563# a_751_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X4 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X5 a_446_3055# MODE_VCCHIB_LV_N VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X6 VCCHIB a_446_3055# OUT_N VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.25
X7 VSSD a_446_3055# OUT_N VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X8 a_751_595# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.8
X9 a_751_595# a_591_563# a_538_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.8
X10 VSSD OUT_N OUT VSSD sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X11 VCCHIB MODE_VCCHIB_LV_N a_612_3332# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.25
X12 VSSD MODE_VCCHIB_LV_N a_446_3055# VSSD sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X13 a_446_3055# a_591_563# a_612_3332# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X14 a_612_3332# a_591_563# a_446_3055# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X15 a_446_3055# a_591_563# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X16 a_751_595# a_591_563# a_538_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.8
X17 VSSD OUT_N OUT VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X18 VSSD IN_H a_751_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X19 a_751_595# IN_H a_591_563# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X20 a_591_563# IN_H a_612_2476# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.8
X21 a_591_563# IN_H a_751_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.8
X22 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0 ps=0 w=5 l=0.8
X23 a_538_595# MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.25
X24 a_612_2476# IN_H a_591_563# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.8
X25 VSSD a_591_563# a_446_3055# VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X26 OUT OUT_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.25
X27 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=0.8
.ends

.subckt sky130_fd_io__gpiov2_in_buf OUT OUT_N MODE_NORMAL_N IN_H IN_VT VTRIP_SEL_H
+ VTRIP_SEL_H_N VDDIO_Q VSSD m1_n467_n748#
X0 a_249_n802# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X1 a_2073_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X2 VSSD a_36_n802# a_2651_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X3 VDDIO_Q VDDIO_Q VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0 ps=0 w=5 l=0.8
X4 a_249_n802# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X5 VDDIO_Q MODE_NORMAL_N a_219_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X6 a_219_1865# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X7 a_249_n802# IN_H a_36_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X8 a_3531_2403# MODE_NORMAL_N a_3358_2403# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X9 a_36_n802# IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X10 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0 ps=0 w=5 l=0.8
X11 a_3358_2403# MODE_NORMAL_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X12 a_2385_1865# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X13 a_36_n802# IN_H a_219_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.8
X14 VDDIO_Q MODE_NORMAL_N a_2073_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X15 VDDIO_Q VTRIP_SEL_H a_3531_2403# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X16 a_249_n802# a_36_n802# a_2073_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.8
X17 VSSD VTRIP_SEL_H a_3358_2403# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X18 VSSD IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X19 a_917_1865# a_973_1767# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X20 VDDIO_Q a_2651_1865# OUT_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X21 OUT OUT_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X22 VSSD IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X23 a_973_1767# a_3358_2403# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X24 a_2651_1865# a_36_n802# a_2385_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X25 VDDIO_Q a_973_1767# a_1761_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X26 a_2073_1865# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X27 a_973_1767# a_3358_2403# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X28 a_249_n802# IN_H a_36_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X29 a_2651_1865# MODE_NORMAL_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X30 a_249_n802# IN_H a_36_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.8
X31 a_36_n802# IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X32 a_1761_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X33 a_2073_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.8
X34 a_249_n802# a_36_n802# a_2073_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X35 a_249_n802# a_36_n802# a_1761_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.8
X36 a_249_n802# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X37 a_3531_2403# MODE_NORMAL_N a_3358_2403# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X38 VSSD IN_VT a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X39 VSSD IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=1.325 ps=10.53 w=5 l=0.8
X40 VSSD VTRIP_SEL_H_N IN_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=1
X41 VDDIO_Q VTRIP_SEL_H a_3531_2403# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X42 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0 ps=0 w=5 l=0.8
X43 VDDIO_Q a_973_1767# a_917_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X44 a_249_n802# a_36_n802# a_1761_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X45 a_917_1865# IN_H a_36_n802# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X46 a_973_1767# a_3358_2403# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X47 a_1761_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X48 a_2651_1865# a_36_n802# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X49 VSSD a_2651_1865# OUT_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X50 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X51 a_1761_1865# a_973_1767# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X52 VSSD MODE_NORMAL_N a_2651_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_ipath_lvls IN_VCCHIB IN_VDDIO MODE_NORMAL_LV MODE_NORMAL_LV_N
+ MODE_VCCHIB_LV MODE_VCCHIB_LV_N VCCHIB VSSD OUT OUT_B a_323_2354#
X0 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X1 VCCHIB MODE_NORMAL_LV_N a_436_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X2 VCCHIB MODE_VCCHIB_LV_N a_1504_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X3 a_823_n317# MODE_NORMAL_LV VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X4 a_114_2354# IN_VDDIO VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X5 a_1679_n317# IN_VCCHIB OUT_B VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X6 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X7 a_1504_2754# IN_VCCHIB OUT_B VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X8 a_323_2354# a_114_2354# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X9 a_436_2754# MODE_NORMAL_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X10 OUT_B a_323_2354# a_436_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X11 VCCHIB OUT_B OUT VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X12 VCCHIB MODE_NORMAL_LV a_114_2354# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.25
X13 VCCHIB OUT_B OUT VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X14 a_823_n317# a_323_2354# OUT_B VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X15 a_1679_n317# MODE_VCCHIB_LV VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X16 a_2141_2754# MODE_NORMAL_LV OUT_B VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X17 a_1504_2754# MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X18 VSSD MODE_NORMAL_LV a_823_n317# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X19 a_316_n17# IN_VDDIO a_114_2354# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.3975 ps=3.53 w=1.5 l=0.5
X20 VSSD MODE_VCCHIB_LV a_1679_n317# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X21 VCCHIB MODE_VCCHIB_LV a_2141_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X22 VCCHIB IN_VDDIO a_114_2354# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X23 OUT_B IN_VCCHIB a_1504_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X24 VSSD MODE_NORMAL_LV a_316_n17# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X25 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X26 a_436_2754# a_323_2354# OUT_B VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X27 a_323_2354# a_114_2354# VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.25
X28 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X29 OUT_B a_323_2354# a_823_n317# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X30 OUT_B IN_VCCHIB a_1679_n317# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
.ends

.subckt sky130_fd_io__gpiov2_inbuf_lvinv_x1 IN VGND VPWR OUT
X0 VPWR IN OUT VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.25
X1 VGND IN OUT VGND sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
.ends

.subckt sky130_fd_io__gpiov2_ibuf_se VTRIP_SEL_H_N VCCHIB ENABLE_VDDIO_LV MODE_NORMAL_N
+ IBUFMUX_OUT IN_VT IN_H VTRIP_SEL_H MODE_VCCHIB_N IBUFMUX_OUT_H sky130_fd_io__gpiov2_in_buf_0/m1_n467_n748#
+ VDDIO_Q VSSD sky130_fd_io__gpiov2_ipath_lvls_0/a_323_2354#
Xsky130_fd_io__gpiov2_ipath_hvls_0 IBUFMUX_OUT_H sky130_fd_io__gpiov2_ipath_hvls_0/OUT_B
+ MODE_NORMAL_N sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT_N
+ sky130_fd_io__gpiov2_in_buf_0/OUT MODE_VCCHIB_N sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL
+ sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB VDDIO_Q VSSD sky130_fd_io__gpiov2_ipath_hvls
Xsky130_fd_io__gpiov2_vcchib_in_buf_0 IN_H sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN
+ VCCHIB VSSD sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT_N
+ sky130_fd_io__gpiov2_vcchib_in_buf
Xsky130_fd_io__gpiov2_in_buf_0 sky130_fd_io__gpiov2_in_buf_0/OUT sky130_fd_io__gpiov2_in_buf_0/OUT_N
+ MODE_NORMAL_N IN_H IN_VT VTRIP_SEL_H VTRIP_SEL_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_in_buf_0/m1_n467_n748#
+ sky130_fd_io__gpiov2_in_buf
Xsky130_fd_io__gpiov2_ipath_lvls_0 sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT sky130_fd_io__gpiov2_in_buf_0/OUT
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN
+ VCCHIB VSSD IBUFMUX_OUT sky130_fd_io__gpiov2_ipath_lvls_0/OUT_B sky130_fd_io__gpiov2_ipath_lvls_0/a_323_2354#
+ sky130_fd_io__gpiov2_ipath_lvls
Xsky130_fd_io__gpiov2_inbuf_lvinv_x1_0 sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN VSSD
+ VCCHIB sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1
Xsky130_fd_io__gpiov2_inbuf_lvinv_x1_1 sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN VSSD
+ VCCHIB sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1
X0 VCCHIB ENABLE_VDDIO_LV sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 VCCHIB sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X2 VSSD MODE_NORMAL_N sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X3 sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X4 sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN ENABLE_VDDIO_LV VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X5 sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB MODE_VCCHIB_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X6 VDDIO_Q MODE_NORMAL_N sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X7 VCCHIB ENABLE_VDDIO_LV sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X8 VCCHIB sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X9 sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X10 sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X11 sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN ENABLE_VDDIO_LV VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X12 VDDIO_Q MODE_NORMAL_N sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X13 sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X14 VSSD ENABLE_VDDIO_LV a_10411_1726# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X15 sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/IN sky130_fd_io__gpiov2_ipath_hvls_0/MODE_NORMAL a_10763_1726# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X16 a_10411_1726# sky130_fd_io__gpiov2_ipath_hvls_0/MODE_VCCHIB sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/IN VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X17 a_10763_1726# ENABLE_VDDIO_LV VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
.ends

.subckt sky130_fd_io__signal_5_sym_hv_local_5term GATE NWELLRING VGND NBODY IN m1_204_67#
X0 IN GATE VGND NBODY sky130_fd_pr__esd_nfet_g5v0d10v5 ad=3.807 pd=12.21 as=3.807 ps=12.21 w=5.4 l=0.6
R0 NBODY m1_534_67# sky130_fd_pr__res_generic_m1 w=0.02 l=5m
R1 NWELLRING m1_204_67# sky130_fd_pr__res_generic_m1 w=0.02 l=5m
.ends

.subckt sky130_fd_io__gpiov2_buf_localesd VTRIP_SEL_H OUT_VT VDDIO_Q VSSD OUT_H IN_H
Xsky130_fd_io__signal_5_sym_hv_local_5term_0 VSSD VDDIO_Q VSSD VSSD OUT_H VDDIO_Q
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_1 VSSD VDDIO_Q OUT_H VSSD VDDIO_Q VDDIO_Q
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__res250only_small_0 IN_H OUT_H sky130_fd_io__res250only_small
X0 OUT_H VTRIP_SEL_H OUT_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=1
.ends

.subckt sky130_fd_io__gpiov2_ipath ENABLE_VDDIO_LV OUT_H VCCHIB DM_H_N[1] DM_H_N[0]
+ DM_H_N[2] INP_DIS_H_N IB_MODE_SEL_H IB_MODE_SEL_H_N VTRIP_SEL_H_N PAD OUT VSSD MODE_VCCHIB_N
+ m1_2058_35701# VDDIO_Q
Xsky130_fd_io__gpiov2_ibuf_se_0 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H_N VCCHIB
+ ENABLE_VDDIO_LV sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N OUT sky130_fd_io__gpiov2_ibuf_se_0/IN_VT
+ sky130_fd_io__gpiov2_ibuf_se_0/IN_H sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H MODE_VCCHIB_N
+ OUT_H PAD VDDIO_Q VSSD m2_15184_37210# sky130_fd_io__gpiov2_ibuf_se
Xsky130_fd_io__gpiov2_buf_localesd_0 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/IN_VT
+ VDDIO_Q VSSD sky130_fd_io__gpiov2_ibuf_se_0/IN_H PAD sky130_fd_io__gpiov2_buf_localesd
X0 a_10749_140# a_11211_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X1 VSSD a_9920_140# a_9864_832# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X2 VSSD DM_H_N[2] a_11331_832# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X3 a_11331_832# a_11211_140# a_10749_140# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X4 VDDIO_Q sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X5 a_9399_166# VTRIP_SEL_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X6 a_10573_140# a_10749_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X7 VDDIO_Q a_10573_140# a_9920_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X8 a_11211_140# a_11563_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X9 VSSD a_10573_140# a_9920_140# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X10 a_11211_140# a_11563_140# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X11 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N a_9399_166# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X12 VDDIO_Q INP_DIS_H_N a_10573_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X13 MODE_VCCHIB_N a_9920_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X14 a_9399_166# VTRIP_SEL_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X15 a_10573_140# a_10749_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X16 VDDIO_Q sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X17 VSSD sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X18 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H VTRIP_SEL_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X19 a_10869_832# a_10749_140# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X20 sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N IB_MODE_SEL_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X21 VDDIO_Q DM_H_N[1] a_11563_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X22 VDDIO_Q IB_MODE_SEL_H MODE_VCCHIB_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X23 a_11563_140# DM_H_N[0] VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X24 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N a_9399_166# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X25 VDDIO_Q INP_DIS_H_N a_10573_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X26 VSSD sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.196 pd=1.96 as=0.098 ps=0.98 w=0.7 l=0.6
X27 a_10573_140# INP_DIS_H_N a_10869_832# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X28 VDDIO_Q a_9920_140# sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X29 VDDIO_Q DM_H_N[2] a_10749_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X30 MODE_VCCHIB_N a_9920_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X31 a_10749_140# a_11211_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X32 a_10216_832# a_9920_140# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X33 sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N IB_MODE_SEL_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X34 VDDIO_Q DM_H_N[1] a_11563_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X35 a_9864_832# IB_MODE_SEL_H_N sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X36 VDDIO_Q a_10573_140# a_9920_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X37 VSSD DM_H_N[1] a_11969_832# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X38 VDDIO_Q IB_MODE_SEL_H MODE_VCCHIB_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X39 a_11563_140# DM_H_N[0] VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X40 a_11211_140# a_11563_140# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X41 MODE_VCCHIB_N IB_MODE_SEL_H a_10216_832# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X42 a_11969_832# DM_H_N[0] a_11563_140# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X43 VDDIO_Q a_9920_140# sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X44 VDDIO_Q DM_H_N[2] a_10749_140# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
.ends

.subckt sky130_fd_io__com_ctl_ls_en_1_v2 DM[1] VCC_IO VPB OUT_H_N OUT_H RST_H SET_H
+ VPWR HLD_H_N a_1150_n777# w_1114_n948# a_1762_n1276# a_n17_1379#
X0 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X7 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X9 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 a_1150_n777# DM[1] a_992_934# w_1114_n948# sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X17 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=1
X18 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X20 a_634_829# a_992_934# a_1150_n777# w_1114_n948# sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X21 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X22 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X23 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X24 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X25 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X26 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X27 a_1762_n1276# DM[1] a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X28 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X29 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X31 a_634_829# a_992_934# a_1762_n1276# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
.ends

.subckt sky130_fd_io__com_ctl_ls_v2 VCC_IO VPB OUT_H_N OUT_H IN RST_H SET_H VPWR HLD_H_N
+ a_n17_1379#
X0 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_634_829# a_992_934# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X7 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X8 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X17 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=1
X18 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 VPWR IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X20 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X22 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X23 a_n17_1379# IN a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X24 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X26 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X27 a_634_829# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X28 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X29 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X31 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
.ends

.subckt sky130_fd_io__com_ctl_lsv2 SET_H HLD_H_N VGND OUT_H OUT_H_N RST_H VPWR VCC_IO
+ m1_5675_1428# w_5775_333# w_4727_n1281# m1_5585_1428# IN
X0 OUT_H a_4739_1530# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X1 OUT_H_N a_4793_n866# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X2 a_4700_638# VPWR a_4933_638# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X3 VGND SET_H a_4739_1530# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X4 VGND a_4739_1530# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X5 VCC_IO a_4793_n866# a_4739_1530# w_4727_n1281# sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X6 a_4700_968# VPWR a_4933_968# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X7 a_4933_968# a_4944_2840# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_4793_n866# RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X9 VGND IN a_4944_2496# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X10 a_4933_968# a_4944_2840# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_4933_638# VPWR a_4700_638# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X12 a_4933_638# HLD_H_N a_4793_n866# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X13 a_4933_968# VPWR a_4700_968# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X14 a_4700_968# VPWR a_4933_968# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X15 VCC_IO a_4793_n866# OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X16 VGND a_4944_2840# a_4933_968# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X17 VGND a_4944_2496# a_4700_638# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VGND a_4944_2496# a_4700_638# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_4933_638# VPWR a_4700_638# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X20 VCC_IO a_4739_1530# a_4793_n866# w_4727_n1281# sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X21 a_4739_1530# a_4793_n866# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=1
X22 a_4944_2840# a_4944_2496# VPWR w_5775_333# sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X23 a_4933_638# VPWR a_4700_638# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X24 a_4944_2840# a_4944_2496# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X25 VGND a_4944_2840# a_4933_968# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X26 a_4793_n866# a_4739_1530# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=1
X27 a_4933_968# VPWR a_4700_968# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X28 VPWR IN a_4944_2496# w_5775_333# sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X29 a_4700_638# a_4944_2496# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X30 a_4700_638# a_4944_2496# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X31 a_4739_1530# HLD_H_N a_4700_968# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
.ends

.subckt sky130_fd_io__com_ctl_ls_1v2 VCC_IO VPB OUT_H_N OUT_H IN RST_H SET_H VPWR
+ HLD_H_N a_n17_1379#
X0 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_634_829# a_992_934# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X7 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X8 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X17 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=1
X18 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 VPWR IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X20 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X22 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X23 a_n17_1379# IN a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X24 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X26 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X27 a_634_829# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X28 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X29 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X31 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_ctl_lsbank VTRIP_SEL_H VTRIP_SEL INP_DIS INP_DIS_H DM[0]
+ DM_H[0] DM_H[2] DM_H_N[2] HLD_I_H_N VCC_IO STARTUP_ST_H STARTUP_RST_H OD_I_H IB_MODE_SEL_H_N
+ sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276# sky130_fd_io__com_ctl_lsv2_0/VCC_IO
+ DM_H[1] INP_DIS_H_N w_15552_2653# m1_2266_545# DM_H_N[1] DM[1] DM_H_N[0] VTRIP_SEL_H_N
+ IB_MODE_SEL VGND IB_MODE_SEL_H VPWR DM[2]
Xsky130_fd_io__com_ctl_ls_en_1_v2_0 DM[1] VCC_IO VPWR DM_H_N[1] DM_H[1] sky130_fd_io__com_ctl_ls_en_1_v2_0/RST_H
+ sky130_fd_io__com_ctl_ls_en_1_v2_0/SET_H VPWR HLD_I_H_N VPWR VPWR sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
+ VGND sky130_fd_io__com_ctl_ls_en_1_v2
Xsky130_fd_io__com_ctl_ls_v2_0 VCC_IO VPWR DM_H_N[2] DM_H[2] DM[2] sky130_fd_io__com_ctl_ls_v2_0/RST_H
+ sky130_fd_io__com_ctl_ls_v2_0/SET_H VPWR HLD_I_H_N VGND sky130_fd_io__com_ctl_ls_v2
Xsky130_fd_io__com_ctl_ls_v2_1 VCC_IO VPWR INP_DIS_H_N INP_DIS_H INP_DIS sky130_fd_io__com_ctl_ls_v2_1/RST_H
+ sky130_fd_io__com_ctl_ls_v2_1/SET_H VPWR HLD_I_H_N VGND sky130_fd_io__com_ctl_ls_v2
Xsky130_fd_io__com_ctl_ls_v2_2 VCC_IO VPWR DM_H_N[0] DM_H[0] DM[0] sky130_fd_io__com_ctl_ls_v2_2/RST_H
+ sky130_fd_io__com_ctl_ls_v2_2/SET_H VPWR HLD_I_H_N VGND sky130_fd_io__com_ctl_ls_v2
Xsky130_fd_io__com_ctl_lsv2_0 sky130_fd_io__com_ctl_lsv2_0/SET_H HLD_I_H_N VGND IB_MODE_SEL_H
+ IB_MODE_SEL_H_N sky130_fd_io__com_ctl_lsv2_0/RST_H VPWR sky130_fd_io__com_ctl_lsv2_0/VCC_IO
+ VGND VPWR w_15552_2653# VGND IB_MODE_SEL sky130_fd_io__com_ctl_lsv2
Xsky130_fd_io__com_ctl_ls_1v2_0 VCC_IO VPWR VTRIP_SEL_H_N VTRIP_SEL_H VTRIP_SEL sky130_fd_io__com_ctl_ls_1v2_0/RST_H
+ sky130_fd_io__com_ctl_ls_1v2_0/SET_H VPWR HLD_I_H_N VGND sky130_fd_io__com_ctl_ls_1v2
R0 m1_5875_412# sky130_fd_io__com_ctl_ls_v2_2/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R1 m1_6420_507# sky130_fd_io__com_ctl_ls_v2_1/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R2 sky130_fd_io__com_ctl_ls_en_1_v2_0/SET_H m1_2266_320# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R3 m1_14183_362# sky130_fd_io__com_ctl_ls_1v2_0/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R4 m2_15089_329# sky130_fd_io__com_ctl_lsv2_0/SET_H sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R5 m1_6620_334# STARTUP_ST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R6 STARTUP_RST_H m1_6420_507# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R7 m1_5875_412# STARTUP_RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R8 m1_6148_320# STARTUP_ST_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R9 m1_10303_506# sky130_fd_io__com_ctl_ls_v2_0/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R10 sky130_fd_io__com_ctl_ls_v2_1/RST_H m1_6620_334# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R11 m1_14183_362# OD_I_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R12 sky130_fd_io__com_ctl_ls_v2_2/SET_H m1_6148_320# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R13 OD_I_H m1_10303_543# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R14 m1_10029_412# OD_I_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R15 m2_15027_104# sky130_fd_io__com_ctl_lsv2_0/SET_H sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R16 m1_6707_412# sky130_fd_io__com_ctl_ls_v2_1/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R17 m1_6421_319# STARTUP_ST_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R18 m2_14799_410# OD_I_H sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R19 m1_14456_624# sky130_fd_io__com_ctl_ls_1v2_0/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R20 m1_5955_333# STARTUP_ST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R21 m1_14457_430# OD_I_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R22 sky130_fd_io__com_ctl_ls_v2_1/SET_H m1_6421_356# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R23 m2_14799_410# sky130_fd_io__com_ctl_lsv2_0/RST_H sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R24 VGND m2_15089_329# sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R25 VGND m1_14456_624# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R26 sky130_fd_io__com_ctl_ls_v2_2/RST_H m1_5955_370# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R27 sky130_fd_io__com_ctl_ls_1v2_0/SET_H m1_14457_467# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R28 m1_10109_333# VGND sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R29 m1_10302_320# VGND sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R30 m1_2553_412# m1_2266_545# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R31 m1_2267_506# sky130_fd_io__com_ctl_ls_en_1_v2_0/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R32 sky130_fd_io__com_ctl_ls_v2_0/RST_H m1_10109_370# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R33 sky130_fd_io__com_ctl_ls_v2_0/SET_H m1_10302_320# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R34 m1_2266_545# m1_2267_543# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R35 m1_14263_617# sky130_fd_io__com_ctl_ls_1v2_0/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R36 m1_2467_333# VGND sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R37 VGND m1_14263_654# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R38 sky130_fd_io__com_ctl_ls_en_1_v2_0/RST_H m1_2467_370# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R39 m1_6149_506# sky130_fd_io__com_ctl_ls_v2_2/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R40 m1_14911_509# sky130_fd_io__com_ctl_lsv2_0/RST_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R41 m2_14990_104# OD_I_H sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R42 m1_10029_412# sky130_fd_io__com_ctl_ls_v2_0/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R43 STARTUP_RST_H m1_6149_543# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R44 m1_2553_412# sky130_fd_io__com_ctl_ls_en_1_v2_0/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R45 VGND m1_14911_546# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R46 m1_2266_320# VGND sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R47 m1_6744_412# STARTUP_RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
.ends

.subckt sky130_fd_io__com_ctl_ls set_h rst_h hld_h_n in out_h vpwr vcc_io vpb out_h_n
+ a_n17_1379#
X0 a_361_1391# vpwr a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 vcc_io a_130_181# out_h vcc_io sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# vpwr a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# hld_h_n a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_634_829# a_992_934# vpwr vpb sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X7 a_361_1391# vpwr a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X8 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 out_h_n a_65_861# vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# hld_h_n a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 out_h a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X17 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=1
X18 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 vpwr in a_992_934# vpb sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X20 a_957_1391# vpwr a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# a_65_861# out_h_n a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X22 a_130_181# a_65_861# vcc_io vcc_io sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X23 a_n17_1379# in a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X24 a_724_1391# vpwr a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X26 a_957_1391# vpwr a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X27 a_634_829# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X28 a_130_181# set_h a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X29 a_724_1391# vpwr a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_128_1391# vpwr a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X31 a_n17_1379# rst_h a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
.ends

.subckt sky130_fd_io__com_ctl_hldv2 HLD_OVR VCC_IO VGND HLD_I_H_N OD_I_H HLD_I_H a_8218_3918#
+ a_3023_3554# m2_3556_4143# m1_3684_4201# a_2671_3554# m2_3665_4182# VPWR
Xsky130_fd_io__com_ctl_ls_0 VGND sky130_fd_io__com_ctl_ls_0/rst_h sky130_fd_io__com_ctl_ls_0/hld_h_n
+ HLD_OVR sky130_fd_io__com_ctl_ls_0/out_h VPWR VCC_IO VPWR sky130_fd_io__com_ctl_ls_0/out_h_n
+ VGND sky130_fd_io__com_ctl_ls
X0 VCC_IO sky130_fd_io__com_ctl_ls_0/hld_h_n a_3743_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 VGND a_3743_3580# a_4447_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X2 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X3 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X4 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X5 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X6 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X7 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X8 VCC_IO sky130_fd_io__com_ctl_ls_0/rst_h a_7214_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X9 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X10 OD_I_H a_7214_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X11 VCC_IO a_7214_3580# OD_I_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X12 VCC_IO OD_I_H a_8391_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X13 VGND a_2671_3554# sky130_fd_io__com_ctl_ls_0/rst_h VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X14 VCC_IO a_3023_3554# a_2967_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X15 VGND sky130_fd_io__com_ctl_ls_0/hld_h_n a_3743_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X16 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X17 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X18 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X19 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X20 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X21 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X22 OD_I_H a_7214_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X23 VCC_IO a_7214_3580# OD_I_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X24 a_8391_3918# a_8271_3554# a_8218_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X25 a_8743_3918# sky130_fd_io__com_ctl_ls_0/hld_h_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X26 a_2967_3918# a_2671_3554# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X27 a_3743_3580# sky130_fd_io__com_ctl_ls_0/hld_h_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X28 a_3743_3580# sky130_fd_io__com_ctl_ls_0/hld_h_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X29 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X30 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X31 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X32 a_8271_3554# sky130_fd_io__com_ctl_ls_0/out_h a_8743_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X33 a_5855_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X34 VGND a_3743_3580# a_4447_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X35 VCC_IO a_2671_3554# sky130_fd_io__com_ctl_ls_0/rst_h VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
R0 HLD_I_H a_3743_3580# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X36 a_5855_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X37 VGND sky130_fd_io__com_ctl_ls_0/rst_h a_7214_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X38 sky130_fd_io__com_ctl_ls_0/hld_h_n a_2967_3918# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X39 VCC_IO sky130_fd_io__com_ctl_ls_0/hld_h_n a_3743_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X40 VCC_IO sky130_fd_io__com_ctl_ls_0/hld_h_n a_3743_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X41 VGND a_7214_3580# OD_I_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X42 VGND OD_I_H a_8218_3918# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X43 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X44 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X45 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X46 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X47 OD_I_H a_7214_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X48 a_2967_3918# a_3023_3554# a_2967_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X49 a_4447_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X50 VGND a_3743_3580# a_5855_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X51 VGND a_3743_3580# a_5855_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X52 OD_I_H a_7214_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X53 a_3743_3580# sky130_fd_io__com_ctl_ls_0/hld_h_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X54 a_8218_3918# a_8271_3554# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X55 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X56 a_8271_3554# sky130_fd_io__com_ctl_ls_0/hld_h_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X57 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X58 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X59 VCC_IO a_7214_3580# OD_I_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X60 a_4447_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X61 VGND a_3743_3580# a_4447_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X62 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X63 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
R1 a_4447_3580# HLD_I_H_N sky130_fd_pr__res_generic_m1 w=0.23 l=0.025
X64 a_2967_3918# a_2671_3554# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X65 a_5855_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X66 VCC_IO sky130_fd_io__com_ctl_ls_0/rst_h a_7214_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
R2 HLD_I_H_N a_5855_3580# sky130_fd_pr__res_generic_m1 w=0.23 l=0.025
X67 a_3743_3580# sky130_fd_io__com_ctl_ls_0/hld_h_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X68 VCC_IO a_7214_3580# OD_I_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X69 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X70 VGND sky130_fd_io__com_ctl_ls_0/out_h a_8271_3554# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.196 pd=1.96 as=0.098 ps=0.98 w=0.7 l=0.6
X71 VCC_IO OD_I_H a_8391_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X72 VCC_IO a_3023_3554# a_2967_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X73 sky130_fd_io__com_ctl_ls_0/hld_h_n a_2967_3918# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.1855 ps=1.93 w=0.7 l=0.6
X74 VGND sky130_fd_io__com_ctl_ls_0/hld_h_n a_3743_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X75 VGND a_3743_3580# a_4447_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X76 a_4447_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X77 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X78 a_5855_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X79 VCC_IO a_2671_3554# sky130_fd_io__com_ctl_ls_0/rst_h VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X80 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X81 VGND a_3743_3580# a_5855_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X82 VCC_IO a_3743_3580# a_5855_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X83 OD_I_H a_7214_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X84 VCC_IO sky130_fd_io__com_ctl_ls_0/hld_h_n a_3743_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X85 OD_I_H a_7214_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X86 a_8391_3918# a_8271_3554# a_8218_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X87 a_8743_3918# sky130_fd_io__com_ctl_ls_0/hld_h_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X88 a_4447_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X89 a_4447_3580# a_3743_3580# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X90 VCC_IO a_3743_3580# a_4447_3580# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X91 a_5855_3580# a_3743_3580# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X92 VGND a_3743_3580# a_5855_3580# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X93 a_3743_3580# sky130_fd_io__com_ctl_ls_0/hld_h_n VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X94 VGND a_7214_3580# OD_I_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X95 a_8271_3554# sky130_fd_io__com_ctl_ls_0/out_h a_8743_3918# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X96 a_2967_3580# a_2671_3554# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X97 sky130_fd_io__com_ctl_ls_0/hld_h_n a_2967_3918# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X98 a_3743_3580# sky130_fd_io__com_ctl_ls_0/hld_h_n VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_ctl DM[0] VTRIP_SEL_H_N DM[2] DM_H[0] DM_H[2] INP_DIS
+ INP_DIS_H_N HLD_OVR VTRIP_SEL VTRIP_SEL_H OD_I_H INP_STARTUP_EN_H IB_MODE_SEL_H_N
+ ENABLE_INP_H HLD_H_N ENABLE_H DM[1] a_11799_3638# li_18199_5031# IB_MODE_SEL_H DM_H_N[0]
+ DM_H_N[1] sky130_fd_io__gpiov2_ctl_lsbank_0/sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
+ DM_H_N[2] DM_H[1] VPWR IB_MODE_SEL HLD_I_H_N HLD_I_OVR_H sky130_fd_io__com_ctl_hldv2_0/HLD_I_H
+ VGND VCC_IO
Xsky130_fd_io__gpiov2_ctl_lsbank_0 VTRIP_SEL_H VTRIP_SEL INP_DIS sky130_fd_io__gpiov2_ctl_lsbank_0/INP_DIS_H
+ DM[0] DM_H[0] DM_H[2] DM_H_N[2] HLD_I_H_N VCC_IO INP_STARTUP_EN_H sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H
+ OD_I_H IB_MODE_SEL_H_N sky130_fd_io__gpiov2_ctl_lsbank_0/sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
+ VCC_IO DM_H[1] INP_DIS_H_N VCC_IO OD_I_H DM_H_N[1] DM[1] DM_H_N[0] VTRIP_SEL_H_N
+ IB_MODE_SEL VGND IB_MODE_SEL_H VPWR DM[2] sky130_fd_io__gpiov2_ctl_lsbank
Xsky130_fd_io__com_ctl_hldv2_0 HLD_OVR VCC_IO VGND HLD_I_H_N OD_I_H sky130_fd_io__com_ctl_hldv2_0/HLD_I_H
+ HLD_I_OVR_H HLD_H_N OD_I_H OD_I_H ENABLE_H OD_I_H VPWR sky130_fd_io__com_ctl_hldv2
X0 INP_STARTUP_EN_H a_11094_4330# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X1 VCC_IO ENABLE_INP_H a_11919_3664# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X2 a_11919_3664# a_11799_3638# sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X3 sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H a_11799_3638# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X4 VCC_IO ENABLE_INP_H a_11919_3664# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X5 a_11094_4330# ENABLE_INP_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X6 VGND ENABLE_INP_H sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X7 VCC_IO OD_I_H a_11094_4330# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X8 INP_STARTUP_EN_H a_11094_4330# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X9 a_11094_4330# ENABLE_INP_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X10 a_11267_4330# ENABLE_INP_H a_11094_4330# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X11 VCC_IO OD_I_H a_11094_4330# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X12 a_11919_3664# a_11799_3638# sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X13 VGND OD_I_H a_11267_4330# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X14 INP_STARTUP_EN_H a_11094_4330# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
.ends

.subckt sky130_fd_io__top_gpiov2 VSSIO_Q PAD_A_NOESD_H ANALOG_POL ENABLE_VDDIO IN_H
+ IN DM[0] DM[1] DM[2] HLD_OVR INP_DIS ENABLE_VDDA_H VTRIP_SEL OE_N OUT SLOW TIE_LO_ESD
+ PAD_A_ESD_0_H ANALOG_SEL ENABLE_INP_H PAD_A_ESD_1_H TIE_HI_ESD ENABLE_H IB_MODE_SEL
+ ENABLE_VSWITCH_H ANALOG_EN sky130_fd_io__overlay_gpiov2_m4_0/sky130_fd_io__top_gpio_pad_0/b_1500_19531#
+ w_9674_16869# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N
+ w_12765_16869# w_12765_14755# w_9674_14653# HLD_H_N VDDIO_Q VSWITCH VSSA PAD VDDIO
+ VCCHIB VDDA AMUXBUS_B AMUXBUS_A VSSIO VCCD VSSD
Xsky130_fd_io__gpio_opathv2_0 sky130_fd_io__gpiov2_ctl_0/HLD_I_OVR_H sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N
+ sky130_fd_io__gpiov2_ctl_0/OD_I_H SLOW VCCD li_3442_6400# li_3302_6400# li_7854_5377#
+ sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpiov2_ctl_0/DM_H[0] sky130_fd_io__gpiov2_ctl_0/DM_H_N[0] li_7943_6398#
+ sky130_fd_io__gpiov2_ctl_0/DM_H[2] sky130_fd_io__gpiov2_ctl_0/DM_H_N[1] VSSD PAD
+ TIE_LO_ESD li_4745_6400# li_7636_6398# sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2]
+ sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H_N li_5278_5352# TIE_HI_ESD VSSD sky130_fd_io__gpiov2_ctl_0/DM_H[1]
+ PAD li_5245_3919# li_9062_7268# sky130_fd_io__gpiov2_ctl_0/DM_H_N[2] li_2678_6400#
+ VDDA li_10974_4971# VCCHIB OE_N OUT VSSD VDDIO sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ li_3958_5352# li_3334_5352# VSSIO sky130_fd_io__gpio_opathv2
Xsky130_fd_io__gpiov2_amux_0 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_13/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_0/ROUT ANALOG_EN ANALOG_POL
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_10/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_10/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_3/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_7/ROUT
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_3/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_13/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_0/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_13/ROUT PAD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N PAD
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ VDDA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_8/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A
+ VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_13/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H PAD VSSA
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_10/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B
+ ANALOG_SEL sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ PAD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N VSSD
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_9/ROUT w_9674_16869# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y
+ AMUXBUS_A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y
+ VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_10/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_6/ROUT
+ VSSA AMUXBUS_B sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/B
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_10/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y
+ sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_3/ROUT sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_6/Y
+ w_12765_16869# VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y
+ w_9674_14653# w_12765_14755# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_3/ROUT
+ VSSD VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_3/ROUT OUT VDDIO_Q
+ PAD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_0/ROUT VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/B
+ VSSD VDDIO_Q VSSD sky130_fd_io__gpiov2_amux
Xsky130_fd_io__res75only_small_0 PAD_A_ESD_1_H sky130_fd_io__res75only_small_1/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_1 sky130_fd_io__res75only_small_1/PAD PAD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_2 PAD_A_ESD_0_H sky130_fd_io__res75only_small_3/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_3 sky130_fd_io__res75only_small_3/PAD PAD sky130_fd_io__res75only_small
Xsky130_fd_io__gpiov2_ipath_0 ENABLE_VDDIO IN_H VCCHIB sky130_fd_io__gpiov2_ctl_0/DM_H_N[1]
+ sky130_fd_io__gpiov2_ctl_0/DM_H_N[0] sky130_fd_io__gpiov2_ctl_0/DM_H_N[2] sky130_fd_io__gpiov2_ctl_0/INP_DIS_H_N
+ sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H_N
+ sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H_N PAD IN VSSD sky130_fd_io__gpiov2_ipath_0/MODE_VCCHIB_N
+ VDDIO VDDIO_Q sky130_fd_io__gpiov2_ipath
Xsky130_fd_io__gpiov2_ctl_0 DM[0] sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H_N DM[2] sky130_fd_io__gpiov2_ctl_0/DM_H[0]
+ sky130_fd_io__gpiov2_ctl_0/DM_H[2] INP_DIS sky130_fd_io__gpiov2_ctl_0/INP_DIS_H_N
+ HLD_OVR VTRIP_SEL sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ctl_0/OD_I_H
+ sky130_fd_io__gpiov2_ctl_0/INP_STARTUP_EN_H sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H_N
+ ENABLE_INP_H HLD_H_N ENABLE_H DM[1] ENABLE_H PAD sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H
+ sky130_fd_io__gpiov2_ctl_0/DM_H_N[0] sky130_fd_io__gpiov2_ctl_0/DM_H_N[1] VSSD sky130_fd_io__gpiov2_ctl_0/DM_H_N[2]
+ sky130_fd_io__gpiov2_ctl_0/DM_H[1] VCCD IB_MODE_SEL sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N
+ sky130_fd_io__gpiov2_ctl_0/HLD_I_OVR_H sky130_fd_io__gpiov2_ctl_0/sky130_fd_io__com_ctl_hldv2_0/HLD_I_H
+ VSSD VDDIO_Q sky130_fd_io__gpiov2_ctl
X0 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT a_2250_17651# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.28 as=4.2 ps=30.56 w=15 l=0.5
X1 a_14092_2778# a_13902_2778# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X2 VCCD a_6895_11435# a_7015_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X3 a_3462_14827# a_3642_14801# a_620_18182# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X4 a_10924_13064# a_334_12102# a_10768_13064# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X5 a_10350_10272# VCCD a_10583_10272# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X6 VSSA a_377_12820# a_2162_14426# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X7 VSSA a_478_17182# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X8 VSSD a_231_9686# a_178_9778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X9 a_9877_11799# a_8765_11461# a_8067_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X10 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H a_1225_12852# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X11 a_10768_13064# a_2250_17651# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X12 a_2159_13760# a_689_12820# a_1024_12357# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X13 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A a_12443_12112# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.15455 pd=1.37 as=0.14 ps=1.28 w=1 l=0.6
X14 a_9406_11799# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X15 VDDA a_184_18182# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X16 VSWITCH a_1024_12357# a_387_12076# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=2
X17 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X18 VDDA a_497_17084# a_229_14828# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=1
X19 a_324_14186# a_689_12820# a_789_14186# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X20 a_620_17850# a_178_9778# a_2080_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X21 a_10406_10767# a_7173_10183# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X22 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N a_184_18182# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X23 w_12765_16869# sky130_fd_io__gpiov2_ctl_0/sky130_fd_io__com_ctl_hldv2_0/HLD_I_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.1176 pd=1.4 as=0.1176 ps=1.4 w=0.42 l=0.5
X24 a_1072_12852# VCCD a_593_13378# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_789_14186# a_689_12820# a_324_14186# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X26 VSSA a_478_17182# a_184_18182# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X27 w_9674_14653# a_6367_11435# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_6/ROUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X28 a_620_18182# a_184_18182# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X29 a_1079_9778# a_282_14802# a_926_9778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X30 a_6367_11435# a_6543_11435# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X31 a_1225_14186# a_689_12820# a_1072_14186# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X32 a_8699_10272# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X33 a_11173_10272# VCCD a_10940_10272# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X34 a_9067_10698# VCCD a_8699_10272# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X35 a_2250_17651# a_7173_10183# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X36 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X37 a_3218_11709# ENABLE_VSWITCH_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X38 a_1077_11842# a_1024_11940# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X39 VSSA VSSA a_387_12076# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X40 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H a_1225_14186# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X41 VSSD a_6895_11435# a_7015_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X42 VDDA ENABLE_VDDA_H a_195_17182# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X43 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A a_11131_11430# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.15455 ps=1.37 w=0.42 l=0.5
X44 a_643_12102# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X45 a_8067_11435# a_8765_11461# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.196 ps=1.96 w=0.7 l=0.6
X46 a_229_14828# a_282_14802# a_382_14828# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X47 VSSD ANALOG_EN a_13816_1289# VSSD sky130_fd_pr__nfet_01v8 ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
R0 PAD PAD_A_NOESD_H sky130_fd_pr__res_generic_m3 w=1.07 l=0.035
X48 a_7367_11461# a_7015_11461# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X49 w_9674_14653# sky130_fd_io__gpiov2_ctl_0/sky130_fd_io__com_ctl_hldv2_0/HLD_I_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.1176 pd=1.4 as=0.1176 ps=1.4 w=0.42 l=0.5
X50 a_593_13760# VCCD a_1072_14186# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X51 a_2982_13760# a_689_12820# a_2162_14426# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X52 a_6895_11435# a_7539_11435# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X53 VSWITCH a_387_12076# a_334_12102# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X54 a_643_12102# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X55 a_14092_2778# VCCD a_14053_2496# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X56 a_7539_11435# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X57 VSWITCH a_1225_12852# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X58 VSSA a_387_12076# a_334_12102# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X59 VSWITCH a_1024_12357# a_2162_14426# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X60 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X61 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_8765_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X62 a_2749_13760# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X63 a_14397_2496# VCCD a_13902_2778# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X64 VCCD a_10643_12610# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.15455 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.5
X65 VSSA a_787_17182# a_2080_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X66 a_9350_10698# VCCD a_8871_10272# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X67 a_6543_11435# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X68 a_13970_2496# a_13760_1103# a_14053_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X69 a_324_14186# a_377_12820# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X70 VSSA a_377_12820# a_324_14186# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X71 a_2080_14827# a_1079_9778# a_184_17734# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X72 VSSD a_7173_10183# a_2250_17651# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X73 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N a_184_18182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X74 VSSA a_195_17182# w_12765_16869# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.1176 pd=1.4 as=0.1176 ps=1.4 w=0.42 l=0.5
X75 a_1072_12852# a_689_12820# a_1225_12852# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X76 a_593_13760# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
R1 PAD_A_NOESD_H PAD sky130_fd_pr__res_generic_m4 w=12.37 l=0.035
X77 VDDIO_Q a_2250_17651# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.28 as=2.1 ps=15.28 w=15 l=0.5
X78 a_2392_13760# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X79 a_178_9778# a_282_14802# a_643_9778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X80 VCCD a_6367_11435# a_6314_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X81 VSSA sky130_fd_io__gpiov2_ctl_0/sky130_fd_io__com_ctl_hldv2_0/HLD_I_H w_9674_16869# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.1176 pd=1.4 as=0.1176 ps=1.4 w=0.42 l=0.5
X82 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H a_231_9686# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X83 a_178_9778# a_1079_9778# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X84 VSWITCH a_1077_11842# a_1024_11940# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=1
X85 a_2159_13760# VCCD a_2392_13760# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X86 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A a_11131_11430# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.15455 pd=1.37 as=0.14 ps=1.28 w=1 l=0.6
X87 a_11523_13190# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X88 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H a_1225_14186# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X89 VSSA a_231_9686# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X90 a_787_17182# a_229_14828# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X91 VSSD a_10643_12610# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.47105 pd=3.65 as=0 ps=0 w=0.42 l=0.5
X92 a_7659_11461# a_7539_11435# a_6895_11435# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X93 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X94 VSSD a_3642_14801# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X95 a_2250_17651# a_7173_10183# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X96 a_421_13760# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X97 VCCD ANALOG_EN a_13816_1289# VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.295 ps=2.59 w=1 l=0.25
X98 VSSA a_195_17182# w_9674_14653# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.1176 pd=1.4 as=0.1176 ps=1.4 w=0.42 l=0.5
X99 a_789_12852# VCCD a_421_13378# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X100 VDDA a_620_18182# a_184_18182# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=1
X101 a_689_12820# a_1024_11940# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X102 VSSA sky130_fd_io__gpiov2_ctl_0/sky130_fd_io__com_ctl_hldv2_0/HLD_I_H w_12765_14755# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.1176 pd=1.4 as=0.1176 ps=1.4 w=0.42 l=0.5
X103 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_178_9778# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X104 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_3642_14801# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X105 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_10705_12172# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X106 a_14397_2496# a_13816_1289# a_13970_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X107 a_10643_12610# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.47105 ps=3.65 w=0.42 l=0.5
X108 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y a_10940_10272# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X109 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y a_7370_13247# VSSD sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X110 a_14053_2496# VCCD a_14092_2778# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X111 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X112 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X113 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y a_7625_13629# VSSD sky130_fd_pr__nfet_01v8 ad=0.2436 pd=1.42 as=0.1008 ps=1.08 w=0.84 l=0.15
X114 VSSD a_6367_11435# a_6314_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
R2 PAD_A_NOESD_H PAD sky130_fd_pr__res_generic_m3 w=12.37 l=0.035
X115 a_1024_12357# a_2162_14426# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X116 a_7621_13247# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y VCCD VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.54 as=0.189 ps=1.56 w=1.26 l=0.15
X117 a_7625_13629# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1008 pd=1.08 as=0.1176 ps=1.12 w=0.84 l=0.15
X118 a_12162_13064# a_334_12102# a_12006_13064# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X119 a_324_14186# a_1225_14186# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X120 VDDA a_497_17084# a_478_17182# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X121 VSSD a_178_9778# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X122 a_2250_17651# a_7173_10183# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X123 a_7621_13247# a_7370_13247# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.3339 pd=3.05 as=0.3591 ps=3.09 w=1.26 l=0.15
X124 a_10705_12172# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_10705_12016# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X125 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H a_1225_12852# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X126 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X127 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X128 a_14053_2496# a_13760_1103# a_13970_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X129 a_10705_11704# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.47105 ps=3.65 w=5 l=0.5
X130 VSSD a_11131_11430# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.47105 pd=3.65 as=0 ps=0 w=0.42 l=0.5
X131 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_8300_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X132 VSSA ENABLE_VSWITCH_H a_342_11805# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.1855 ps=1.93 w=0.7 l=0.6
X133 a_421_13378# VCCD a_789_12852# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X134 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A a_12443_12112# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.47105 pd=3.65 as=0.1113 ps=1.37 w=0.42 l=0.5
X135 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_12897_12172# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X136 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y a_8871_10272# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X137 a_13970_2496# a_13816_1289# a_14397_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X138 VCCD a_6895_11435# a_7015_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X139 a_8699_10272# VCCD a_9067_10698# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X140 a_620_17850# a_184_17734# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X141 VSSD a_7173_10183# a_2250_17651# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X142 a_9877_11799# a_8765_11461# a_8067_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X143 VSSD a_7173_10183# a_2250_17651# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X144 a_2250_17651# a_7173_10183# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X145 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT a_2250_17651# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=4.2 pd=30.56 as=2.1 ps=15.28 w=15 l=0.5
X146 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H a_1225_12852# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X147 a_14397_2496# a_13816_1289# a_13970_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X148 VSSD sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N a_13970_2496# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X149 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X150 a_497_17084# a_195_17182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X151 a_2080_14827# a_178_9778# a_620_17850# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X152 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X153 a_447_9352# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X154 a_2080_14827# a_1079_9778# a_184_17734# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X155 a_7173_10183# a_231_9686# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X156 a_9406_11799# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X157 a_12897_12172# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_12897_12016# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X158 a_620_17850# a_178_9778# a_2080_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X159 a_1072_14186# VCCD a_593_13760# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X160 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A a_12443_12112# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.15455 ps=1.37 w=0.42 l=0.5
X161 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A a_8699_10272# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X162 VDDIO_Q a_3642_14801# a_4110_14801# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X163 a_12897_11704# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.47105 ps=3.65 w=5 l=0.5
X164 VCCD a_8067_11435# a_6543_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X165 VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y a_593_13378# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X166 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT a_2250_17651# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.28 as=2.1 ps=15.28 w=15 l=0.5
X167 a_447_9352# VCCD a_926_9778# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X168 a_497_17084# a_231_9686# a_382_14828# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X169 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_8473_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X170 VDDIO_Q a_2250_17651# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.28 as=2.1 ps=15.28 w=15 l=0.5
X171 VCCD a_6543_11435# a_6367_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X172 w_9674_16869# a_195_17182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.1176 pd=1.4 as=0.1176 ps=1.4 w=0.42 l=0.5
X173 a_3642_14801# a_282_14802# a_9067_10698# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X174 VSSA a_1225_12852# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X175 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A a_11523_13190# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.15455 ps=1.37 w=0.42 l=0.5
X176 a_13970_2496# a_13816_1289# a_14397_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X177 a_643_9778# a_282_14802# a_178_9778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X178 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H a_1225_14186# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X179 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y a_447_9352# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X180 a_13902_2778# VCCD a_14397_2496# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X181 VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A a_421_13378# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X182 a_195_17182# ENABLE_VDDA_H VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X183 a_14053_2496# a_13760_1103# a_13970_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X184 a_6895_11435# a_7539_11435# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X185 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_11/Y a_7453_13247# VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.189 pd=1.56 as=0.1512 ps=1.5 w=1.26 l=0.15
X186 VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_0/Y a_2749_13760# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X187 a_10643_12610# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.15455 ps=1.37 w=1 l=0.6
X188 a_275_9352# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X189 a_7453_13247# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y a_7370_13247# VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.1512 pd=1.5 as=0.3339 ps=3.05 w=1.26 l=0.15
X190 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H a_9877_11799# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X191 VSSA a_1225_14186# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X192 a_7173_10183# a_282_14802# a_11173_10272# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X193 w_12765_14755# a_195_17182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.1176 pd=1.4 as=0.1176 ps=1.4 w=0.42 l=0.5
X194 a_324_12852# a_689_12820# a_789_12852# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X195 a_787_17182# a_229_14828# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X196 a_184_17734# a_1079_9778# a_2080_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X197 a_6543_11435# a_8067_11435# a_8011_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X198 a_387_12076# a_1024_12357# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=2
X199 a_11173_10272# a_282_14802# a_7173_10183# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X200 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X201 a_10406_10767# a_282_14802# a_10350_10272# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X202 a_789_12852# a_689_12820# a_324_12852# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X203 VSSA a_497_17084# a_478_17182# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X204 a_926_9778# VCCD a_447_9352# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X205 a_7539_11435# a_8300_11461# a_9406_11799# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X206 a_11850_13064# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.47105 ps=3.65 w=5 l=0.5
X207 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X208 a_1225_12852# a_689_12820# a_1072_12852# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X209 VSSD a_13816_1289# a_13760_1103# VSSD sky130_fd_pr__nfet_01v8 ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X210 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A a_2250_17651# a_12162_13064# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X211 VSWITCH ENABLE_VSWITCH_H a_342_11805# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X212 VSSD a_6543_11435# a_6367_11435# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X213 VCCD a_6367_11435# a_6314_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X214 VSWITCH a_324_14186# a_1225_14186# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X215 VDDA a_620_17850# a_184_17734# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=1
X216 a_13970_2496# a_13760_1103# a_14053_2496# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X217 a_9350_10698# a_282_14802# a_4110_14801# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X218 a_1077_11842# a_342_11805# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X219 a_324_12852# a_1225_12852# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X220 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A a_275_9352# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X221 VDDIO_Q a_13902_2778# a_231_9686# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X222 w_12765_14755# a_6367_11435# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_7/ROUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X223 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H a_1225_14186# VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X224 a_9067_10698# a_282_14802# a_3642_14801# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X225 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X226 a_10940_10272# VCCD a_11173_10272# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X227 a_184_17734# a_478_17182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X228 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y a_10583_10272# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X229 a_8300_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X230 VSSA a_1225_14186# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X231 a_497_17084# a_229_14828# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X232 VSSA a_184_17734# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X233 a_2982_13760# VCCD a_2749_13760# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X234 a_789_14186# VCCD a_421_13760# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X235 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H a_8067_11435# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X236 a_7015_11461# a_6895_11435# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X237 VSWITCH a_1077_11842# a_377_12820# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X238 a_8765_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X239 a_1077_11842# a_231_9686# a_3218_11709# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X240 a_2250_17651# a_7173_10183# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X241 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y a_6895_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X242 a_643_9778# VCCD a_275_9352# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X243 VDDIO_Q a_7173_10183# a_2250_17651# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X244 a_324_12852# a_377_12820# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X245 a_14092_2778# VCCD a_14053_2496# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X246 VSSD a_8300_11461# a_7539_11435# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.196 pd=1.96 as=0.098 ps=0.98 w=0.7 l=0.6
X247 VSSA a_377_12820# a_324_12852# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X248 a_184_18182# a_4110_14801# a_3462_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X249 a_11080_13064# a_6314_11461# a_10924_13064# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X250 a_2162_14426# a_377_12820# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X251 a_10350_10272# a_282_14802# a_10406_10767# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X252 a_13970_2496# sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X253 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A a_10643_12610# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X254 VSSA ENABLE_VDDA_H a_382_14828# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X255 a_3462_14827# a_4110_14801# a_184_18182# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X256 a_3642_14801# a_4110_14801# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X257 a_4110_14801# a_282_14802# a_9350_10698# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X258 VCCD a_13816_1289# a_13760_1103# VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.295 ps=2.59 w=1 l=0.25
X259 a_12443_12112# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X260 a_3642_14801# a_231_9686# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X261 VDDIO_Q a_3642_14801# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X262 a_275_9352# VCCD a_643_9778# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X263 a_8473_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N a_8300_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X264 a_7370_13247# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X265 VDDIO_Q a_178_9778# a_1079_9778# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X266 VSSD a_231_9686# a_3642_14801# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X267 a_6367_11435# a_6543_11435# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X268 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X269 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_8300_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X270 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X271 VSSA a_1024_11940# a_689_12820# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X272 a_10583_10272# VCCD a_10350_10272# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X273 a_7015_11461# a_6895_11435# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X274 a_8938_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N a_8765_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X275 a_421_13760# VCCD a_789_14186# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X276 a_1072_14186# a_689_12820# a_1225_14186# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X277 a_3218_11709# a_231_9686# a_1077_11842# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X278 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y a_7659_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X279 a_178_9778# a_231_9686# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X280 w_12765_16869# a_7015_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_9/ROUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X281 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A a_11131_11430# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.47105 pd=3.65 as=0.1113 ps=1.37 w=0.42 l=0.5
X282 a_497_17084# a_231_9686# a_382_14828# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X283 a_7367_11461# a_7015_11461# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X284 VSSD a_231_9686# a_7173_10183# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X285 a_4259_12681# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X286 VSSD a_12443_12112# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.47105 pd=3.65 as=0 ps=0 w=0.42 l=0.5
X287 a_184_18182# a_4110_14801# a_3462_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X288 a_382_14828# a_282_14802# a_229_14828# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X289 a_593_13378# VCCD a_1072_12852# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X290 a_8871_10272# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X291 VSSA a_1225_12852# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.6
X292 a_2162_14426# a_689_12820# a_2982_13760# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X293 a_8871_10272# VCCD a_9350_10698# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X294 a_926_9778# a_282_14802# a_1079_9778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X295 VDDIO_Q a_178_9778# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X296 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_8765_11461# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X297 a_12006_13064# a_7367_11461# a_11850_13064# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X298 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A a_11080_13064# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.47105 pd=3.65 as=0.7 ps=5.28 w=5 l=0.5
X299 VSSD a_7370_13247# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nand2_1_1/B VSSD sky130_fd_pr__nfet_01v8 ad=0.4788 pd=2.82 as=0.2436 ps=1.42 w=0.84 l=0.15
X300 a_1024_12357# a_689_12820# a_2159_13760# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X301 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X302 VSSD a_11523_13190# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=0.5
X303 a_6543_11435# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X304 a_3462_14827# a_787_17182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X305 a_10705_12016# a_643_12102# a_10705_11860# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X306 a_2250_17651# a_7173_10183# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X307 a_2749_13760# VCCD a_2982_13760# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X308 VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/Y a_593_13760# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X309 VCCD a_8067_11435# a_6543_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X310 VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/Y a_2392_13760# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X311 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X312 a_342_11805# ENABLE_VSWITCH_H VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X313 a_6367_11435# a_6543_11435# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X314 a_387_12076# a_231_9686# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X315 a_13902_2778# a_14092_2778# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X316 VCCD a_6543_11435# a_6367_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X317 VSWITCH a_324_12852# a_1225_12852# VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X318 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N a_178_9778# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.6
X319 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_3642_14801# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X320 a_14397_2496# VCCD a_13902_2778# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X321 VDDIO_Q a_7173_10183# a_2250_17651# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X322 VDDIO_Q a_7173_10183# a_2250_17651# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X323 a_13902_2778# sky130_fd_io__gpiov2_ctl_0/sky130_fd_io__com_ctl_hldv2_0/HLD_I_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X324 a_10705_11860# a_4259_12681# a_10705_11704# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X325 VSWITCH a_1225_12852# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X326 a_593_13378# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/Y VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X327 VSSA sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_9/A a_421_13760# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X328 a_1077_11842# a_231_9686# a_3218_11709# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X329 a_387_12076# a_1024_12357# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X330 VSSD a_14092_2778# a_282_14802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X331 VSSD sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N a_13970_2496# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X332 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A a_11523_13190# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.15455 pd=1.37 as=0.14 ps=1.28 w=1 l=0.6
X333 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A a_11523_13190# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.47105 pd=3.65 as=0.1113 ps=1.37 w=0.42 l=0.5
X334 a_7367_11461# a_7015_11461# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X335 a_13970_2496# sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X336 a_12897_12016# a_643_12102# a_12897_11860# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X337 a_11131_11430# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X338 a_195_17182# ENABLE_VDDA_H VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X339 a_2250_17651# a_7173_10183# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X340 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H a_9877_11799# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X341 a_382_14828# a_282_14802# a_229_14828# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X342 VSSD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N a_8938_11461# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X343 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_8/ROUT a_7015_11461# w_9674_16869# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X344 a_421_13378# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_8/A VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X345 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X346 VSWITCH a_1225_14186# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X347 a_3462_14827# a_3642_14801# a_620_18182# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X348 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X349 VDDIO_Q a_10406_10767# a_7173_10183# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X350 a_8011_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X351 a_620_18182# a_3642_14801# a_3462_14827# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X352 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X353 a_7539_11435# a_8300_11461# a_9406_11799# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X354 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y a_7621_13247# VCCD sky130_fd_pr__pfet_01v8_hvt ad=0.4786 pd=3.44 as=0.1764 ps=1.54 w=1.26 l=0.15
X355 a_282_14802# a_14092_2778# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X356 a_2392_13760# VCCD a_2159_13760# VSSA sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X357 a_12897_11860# a_4259_12681# a_12897_11704# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X358 VSSA a_1077_11842# a_377_12820# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X359 a_2250_17651# a_7173_10183# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.6
X360 VDDA a_184_17734# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X361 a_4259_12681# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.3975 ps=3.53 w=1.5 l=0.5
X362 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT a_2250_17651# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.28 as=2.1 ps=15.28 w=15 l=0.5
X363 a_10940_10272# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_1/Y VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X364 a_3218_11709# a_282_14802# a_1024_11940# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X365 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N a_184_17734# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X366 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_4/ROUT a_387_12076# VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.56 w=5 l=0.5
X367 VDDIO_Q a_2250_17651# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.28 as=2.1 ps=15.28 w=15 l=0.5
X368 a_231_9686# a_13902_2778# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X369 a_8300_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X370 a_1024_11940# a_282_14802# a_3218_11709# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X371 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H a_1225_12852# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.6
X372 a_3218_11709# a_282_14802# a_1024_11940# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X373 VSWITCH a_1225_14186# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X374 a_13902_2778# VCCD a_14397_2496# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X375 VSSIO_Q a_387_12076# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__res75only_small_5/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.56 as=0.7 ps=5.28 w=5 l=0.5
X376 a_14053_2496# VCCD a_14092_2778# VSSD sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X377 a_7015_11461# a_6895_11435# VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X378 a_8765_11461# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N VCCD VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X379 a_382_14828# a_231_9686# a_497_17084# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X380 VCCD sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y a_6895_11435# VCCD sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X381 a_10583_10272# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_5/Y VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X382 sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H a_478_17182# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
.ends

.subckt sky130_ef_io__gpiov2_pad DM[0] IB_MODE_SEL ENABLE_H ENABLE_INP_H SLOW VTRIP_SEL
+ ENABLE_VDDIO ENABLE_VDDA_H PAD_A_NOESD_H ANALOG_POL HLD_H_N w_9674_16462# DM[1]
+ w_12765_14348# DM[2] w_9674_14246# PAD_A_ESD_1_H TIE_HI_ESD ENABLE_VSWITCH_H TIE_LO_ESD
+ OE_N w_12765_16462# AMUXBUS_B ANALOG_SEL VSWITCH AMUXBUS_A IN_H VDDIO INP_DIS OUT
+ HLD_OVR VCCD PAD VCCHIB PAD_A_ESD_0_H ANALOG_EN VSSIO VDDA VDDIO_Q VSSIO_Q VSSA
+ IN VSSD
Xsky130_fd_io__top_gpiov2_0 VSSIO_Q PAD_A_NOESD_H ANALOG_POL ENABLE_VDDIO IN_H IN
+ DM[0] DM[1] DM[2] HLD_OVR INP_DIS ENABLE_VDDA_H VTRIP_SEL OE_N OUT SLOW TIE_LO_ESD
+ PAD_A_ESD_0_H ANALOG_SEL ENABLE_INP_H PAD_A_ESD_1_H TIE_HI_ESD ENABLE_H IB_MODE_SEL
+ ENABLE_VSWITCH_H ANALOG_EN sky130_fd_io__top_gpiov2_0/sky130_fd_io__overlay_gpiov2_m4_0/sky130_fd_io__top_gpio_pad_0/b_1500_19531#
+ w_9674_16462# sky130_fd_io__top_gpiov2_0/sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N
+ w_12765_16462# w_12765_14348# w_9674_14246# HLD_H_N VDDIO_Q VSWITCH VSSA PAD VDDIO
+ VCCHIB VDDA AMUXBUS_B AMUXBUS_A VSSIO VCCD VSSD sky130_fd_io__top_gpiov2
.ends

.subckt sky130_fd_io__sio_clamp_pcap_4x5 a_36_36# a_229_118#
X0 a_36_36# a_229_118# a_36_36# a_36_36# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0 ps=0 w=5 l=4
.ends

.subckt sky130_fd_io__pad_esd m4_960_20017# m5_1354_20500#
R0 m4_960_20017# m5_1354_20500# sky130_fd_pr__res_generic_m5 w=252.96001 l=0.1
.ends

.subckt sky130_fd_io__com_busses_esd sky130_fd_io__com_bus_hookup_0/VCCHIB sky130_fd_io__pad_esd_0/m5_1354_20500#
+ sky130_fd_io__com_bus_hookup_0/VSSD sky130_fd_io__pad_esd_0/m4_960_20017# sky130_fd_io__com_bus_hookup_0/AMUXBUS_A
+ sky130_fd_io__com_bus_hookup_0/VCCD sky130_fd_io__com_bus_hookup_0/AMUXBUS_B sky130_fd_io__com_bus_hookup_0/VDDIO
+ sky130_fd_io__com_bus_hookup_0/VSSA sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_bus_hookup_0/VSWITCH
+ sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_bus_hookup_0/VDDIO_Q sky130_fd_io__com_bus_hookup_0/VSSIO_Q
Xsky130_fd_io__pad_esd_0 sky130_fd_io__pad_esd_0/m4_960_20017# sky130_fd_io__pad_esd_0/m5_1354_20500#
+ sky130_fd_io__pad_esd
.ends

.subckt sky130_fd_io__esd_rcclamp_nfetcap a_179_100# a_n14_18#
X0 a_n14_18# a_179_100# a_n14_18# a_n14_18# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0 ps=0 w=5 l=8
.ends

.subckt sky130_fd_io__top_ground_hvc_wpad VCCHIB VDDA VDDIO_Q VSSIO_Q G_PAD PADISOR
+ PADISOL DRN_HVC SRC_BDY_HVC OGC_HVC G_CORE AMUXBUS_B VSSIO VDDIO VSSD VSWITCH VSSA
+ AMUXBUS_A VCCD
Xsky130_fd_io__sio_clamp_pcap_4x5_0 SRC_BDY_HVC a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__com_busses_esd_0 VCCHIB G_PAD VSSD G_CORE AMUXBUS_A VCCD AMUXBUS_B
+ VDDIO VSSA VSSIO VSWITCH VDDA VDDIO_Q VSSIO_Q sky130_fd_io__com_busses_esd
Xsky130_fd_io__sio_clamp_pcap_4x5_1[0] SRC_BDY_HVC a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__sio_clamp_pcap_4x5_1[1] SRC_BDY_HVC a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__sio_clamp_pcap_4x5_1[2] SRC_BDY_HVC a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|0] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|0] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|0] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|1] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|1] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|1] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|2] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|2] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|2] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|3] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|3] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|3] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|4] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|4] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|4] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
X0 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X1 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X2 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X3 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X4 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.855 ps=14.53 w=7 l=0.5
X5 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X6 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X7 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X8 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X9 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X10 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X11 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X12 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X13 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X14 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X15 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X16 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X17 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X18 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X19 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X20 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X21 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X22 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X23 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X24 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X25 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X26 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X27 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X28 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X29 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X30 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X31 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X32 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X33 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X34 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X35 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X36 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X37 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X38 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X39 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X40 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X41 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X42 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X43 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X44 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X45 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X46 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X47 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X48 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X49 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X50 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X51 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X52 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X53 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X54 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X55 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X56 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X57 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X58 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X59 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X60 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X61 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X62 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X63 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
R0 G_CORE PADISOL sky130_fd_pr__res_generic_m3 w=11.825 l=10m
X64 SRC_BDY_HVC a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0 ps=0 w=5 l=4
X65 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X66 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X67 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X68 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X69 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X70 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X71 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X72 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X73 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X74 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X75 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X76 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X77 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X78 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X79 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X80 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X81 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X82 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X83 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X84 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X85 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X86 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X87 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X88 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X89 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X90 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X91 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X92 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X93 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X94 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X95 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X96 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X97 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X98 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X99 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X100 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
R1 G_CORE PADISOR sky130_fd_pr__res_generic_m3 w=11.825 l=10m
X101 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X102 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X103 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X104 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X105 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X106 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X107 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X108 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X109 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X110 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X111 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X112 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X113 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X114 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X115 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X116 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X117 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X118 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X119 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X120 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X121 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X122 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X123 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X124 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X125 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X126 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X127 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X128 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X129 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X130 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X131 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X132 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X133 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X134 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X135 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X136 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X137 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X138 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X139 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X140 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X141 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X142 DRN_HVC a_214_8638# sky130_fd_pr__res_generic_po w=0.33 l=700
X143 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X144 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X145 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=1.855 pd=14.53 as=0.98 ps=7.28 w=7 l=0.5
X146 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X147 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X148 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X149 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X150 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X151 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.855 ps=14.53 w=7 l=0.5
X152 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X153 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X154 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X155 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X156 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X157 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X158 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X159 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X160 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X161 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X162 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X163 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X164 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X165 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X166 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X167 a_1672_8638# a_214_8638# sky130_fd_pr__res_generic_po w=0.33 l=1.55k
X168 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X169 a_1268_5934# a_1672_8638# sky130_fd_pr__res_generic_po w=0.33 l=470
X170 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X171 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X172 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X173 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X174 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X175 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X176 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X177 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X178 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X179 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X180 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X181 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X182 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X183 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X184 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X185 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X186 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X187 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X188 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X189 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X190 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X191 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X192 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X193 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X194 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X195 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X196 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X197 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X198 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X199 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X200 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X201 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X202 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X203 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X204 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X205 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=1.855 pd=14.53 as=0.98 ps=7.28 w=7 l=0.5
X206 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X207 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X208 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X209 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X210 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
.ends

.subckt sky130_ef_io__vssio_hvc_clamped_pad VDDA VSSD VSSA AMUXBUS_A AMUXBUS_B VSSIO_PAD
+ VDDIO_Q VDDIO VSSIO VSWITCH VSSIO_Q VCCHIB VCCD
Xsky130_fd_io__top_ground_hvc_wpad_2 VCCHIB VDDA VDDIO_Q VSSIO_Q VSSIO_PAD VSSIO_Q
+ VSSIO_Q VDDIO VSSIO VDDIO VSSIO AMUXBUS_B VSSIO VDDIO VSSD VSWITCH VSSA AMUXBUS_A
+ VCCD sky130_fd_io__top_ground_hvc_wpad
.ends

.subckt chip_io_gpio_connects_horiz tie_lo_esd in tie_hi_esd enable_vddio slow pad_a_esd_0_h
+ pad_a_esd_1_h dm[1] pad_a_noesd_h analog_en dm[0] analog_pol inp_dis enable_inp_h
+ enable_h hld_h_n analog_sel dm[2] hld_ovr out enable_vswitch_h enable_vdda_h vtrip_sel
+ ib_mode_sel oe_n in_h one zero constant_block_0/vccd VSUBS
Xconstant_block_0 one constant_block_0/vccd zero VSUBS constant_block
.ends

.subckt sky130_fd_io__hvc_clampv2 m2_5179_0# w_1040_5785# sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20500#
+ m3_10082_12712# m3_103_12712# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q
+ w_2676_441# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO m3_99_0# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD
Xsky130_fd_io__sio_clamp_pcap_4x5_0[0] w_2676_441# a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__sio_clamp_pcap_4x5_0[1] w_2676_441# a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__sio_clamp_pcap_4x5_0[2] w_2676_441# a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__com_busses_esd_0 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20500# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD
+ m3_99_0# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q sky130_fd_io__com_busses_esd
Xsky130_fd_io__sio_clamp_pcap_4x5_1 w_2676_441# a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|0] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|0] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|0] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|1] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|1] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|1] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|2] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|2] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|2] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|3] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|3] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|3] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|4] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|4] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|4] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
X0 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X1 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X2 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X3 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X4 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.855 ps=14.53 w=7 l=0.5
X5 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X6 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X7 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X8 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X9 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X10 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X11 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X12 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X13 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X14 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X15 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X16 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X17 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X18 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X19 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X20 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X21 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X22 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X23 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X24 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X25 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X26 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X27 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X28 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X29 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X30 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X31 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X32 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X33 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X34 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X35 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X36 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X37 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X38 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X39 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X40 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X41 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X42 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X43 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X44 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X45 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X46 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X47 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X48 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X49 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X50 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X51 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X52 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X53 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X54 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X55 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X56 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X57 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X58 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X59 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X60 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X61 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X62 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X63 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X64 w_2676_441# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0 ps=0 w=5 l=4
X65 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X66 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X67 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X68 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X69 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X70 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X71 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X72 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X73 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X74 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X75 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X76 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X77 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X78 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X79 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X80 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X81 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X82 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X83 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X84 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X85 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X86 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X87 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X88 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X89 a_1268_5934# a_1672_8570# sky130_fd_pr__res_generic_po w=0.33 l=470
X90 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X91 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X92 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X93 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X94 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X95 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X96 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X97 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X98 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X99 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X100 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X101 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X102 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X103 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X104 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X105 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X106 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X107 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X108 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X109 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X110 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X111 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X112 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X113 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X114 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X115 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X116 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X117 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X118 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X119 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X120 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X121 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X122 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X123 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X124 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X125 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X126 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X127 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X128 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X129 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X130 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X131 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X132 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X133 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X134 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X135 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X136 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
R0 m3_99_0# m3_103_12712# sky130_fd_pr__res_generic_m3 w=12.125 l=10m
X137 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X138 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X139 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X140 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X141 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X142 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X143 w_1040_5785# a_214_8570# sky130_fd_pr__res_generic_po w=0.33 l=700
X144 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X145 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X146 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=1.855 pd=14.53 as=0.98 ps=7.28 w=7 l=0.5
X147 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X148 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X149 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X150 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X151 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X152 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.855 ps=14.53 w=7 l=0.5
X153 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X154 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X155 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X156 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X157 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X158 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X159 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X160 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X161 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X162 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X163 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X164 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X165 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X166 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X167 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X168 a_1672_8570# a_214_8570# sky130_fd_pr__res_generic_po w=0.33 l=1.55k
X169 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X170 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X171 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X172 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X173 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X174 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X175 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
R1 m3_99_0# m3_10082_12712# sky130_fd_pr__res_generic_m3 w=12.125 l=10m
X176 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X177 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X178 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X179 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X180 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X181 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X182 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X183 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X184 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X185 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X186 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X187 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X188 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X189 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X190 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X191 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X192 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
X193 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X194 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X195 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X196 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X197 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X198 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X199 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X200 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X201 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X202 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X203 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.51 as=6.95 ps=21.39 w=10 l=0.5
X204 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.39 as=15.1 ps=21.51 w=20 l=0.5
X205 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=1.855 pd=14.53 as=0.98 ps=7.28 w=7 l=0.5
X206 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X207 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X208 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X209 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.51 as=13.9 ps=41.39 w=20 l=0.5
X210 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.39 as=7.55 ps=11.51 w=10 l=0.5
.ends

.subckt sky130_fd_io__top_power_hvc_wpadv2 SRC_BDY_HVC OGC_HVC AMUXBUS_B VDDA VSSIO_Q
+ P_PAD PADISOL VDDIO_Q P_CORE PADISOR DRN_HVC VCCHIB VCCD VSWITCH VDDIO VSSA VSSD
+ AMUXBUS_A VSSIO
Xsky130_fd_io__hvc_clampv2_0 OGC_HVC DRN_HVC P_PAD PADISOR PADISOL VDDIO_Q AMUXBUS_B
+ VSSIO_Q SRC_BDY_HVC VCCHIB VSSIO VDDA VDDIO P_CORE VSSD VSWITCH VSSA AMUXBUS_A VCCD
+ sky130_fd_io__hvc_clampv2
.ends

.subckt sky130_ef_io__vddio_hvc_clamped_pad VDDA VSSIO_Q VDDIO VDDIO_Q VSSD VDDIO_PAD
+ VSSA AMUXBUS_B AMUXBUS_A VSWITCH VCCHIB VSSIO VCCD
Xsky130_fd_io__top_power_hvc_wpadv2_2 VSSIO VDDIO AMUXBUS_B VDDA VSSIO_Q VDDIO_PAD
+ VDDIO_Q VDDIO_Q VDDIO VDDIO_Q VDDIO VCCHIB VCCD VSWITCH VDDIO VSSA VSSD AMUXBUS_A
+ VSSIO sky130_fd_io__top_power_hvc_wpadv2
.ends

.subckt sky130_fd_io__gpiovrefv2_res_ladder vrefgen_en_h vrefgen_en_h_n vref<31> vref<30>
+ vref<29> vref<28> vref<27> vref<26> vref<25> vref<24> vref<23> vref<22> vref<21>
+ vref<20> vref<19> vref<18> vref<17> vref<16> vref<15> vref<14> vref<13> vref<12>
+ vref<11> vref<10> vref<9> vref<8> vref<7> vref<6> vref<5> vref<4> vref<3> vref<2>
+ vref<1> vref<0> vssd vddio_q a_9088_3179# a_n252_3179#
X0 vref<31> a_n138_3352# vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X1 vref<14> vref<15> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X2 vref<9> vref<10> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X3 vref<2> vref<3> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X4 vref<24> vref<25> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X5 vref<19> vref<20> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X6 vref<8> vref<9> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X7 vddio_q vrefgen_en_h_n a_n138_3352# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X8 vref<12> vref<13> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X9 vref<7> vref<8> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X10 a_n138_3352# vrefgen_en_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X11 a_12896_38573# a_13320_n869# vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=2.4775k
X12 a_13320_n869# vrefgen_en_h a_11607_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X13 a_11607_n869# vrefgen_en_h a_13320_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X14 vssd vrefgen_en_h a_11607_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X15 vref<6> vref<7> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X16 vssd vrefgen_en_h a_11607_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X17 a_11607_n869# vrefgen_en_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X18 a_13320_n869# vrefgen_en_h a_11607_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X19 a_11607_n869# vrefgen_en_h a_13320_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X20 vref<1> vref<2> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X21 vddio_q vrefgen_en_h_n a_n138_3352# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X22 a_n138_3352# vrefgen_en_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X23 vref<29> vref<30> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X24 a_12896_38573# vref<0> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=2.4775k
X25 vddio_q vrefgen_en_h_n a_n138_3352# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X26 vref<23> vref<24> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X27 a_11607_n869# vrefgen_en_h a_13320_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X28 a_13320_n869# vrefgen_en_h a_11607_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X29 vref<0> vref<1> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X30 vssd vrefgen_en_h a_11607_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X31 a_11607_n869# vrefgen_en_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X32 vref<27> vref<28> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X33 a_11607_n869# vrefgen_en_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X34 vref<5> vref<6> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X35 vref<15> vref<16> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X36 vref<10> vref<11> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X37 vref<28> vref<29> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X38 vref<4> vref<5> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X39 a_13320_n869# vrefgen_en_h a_11607_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X40 a_11607_n869# vrefgen_en_h a_13320_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X41 vref<18> vref<19> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X42 a_n138_3352# vrefgen_en_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X43 a_11607_n869# vrefgen_en_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X44 vssd vrefgen_en_h a_11607_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X45 a_11607_n869# vrefgen_en_h vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X46 vref<22> vref<23> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X47 vref<17> vref<18> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X48 vref<13> vref<14> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X49 vref<26> vref<27> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X50 vref<11> vref<12> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X51 a_n138_3352# vrefgen_en_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X52 vref<21> vref<22> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X53 vref<16> vref<17> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X54 vddio_q vrefgen_en_h_n a_n138_3352# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X55 vref<3> vref<4> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X56 a_n138_3352# vrefgen_en_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X57 vref<30> vref<31> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X58 vref<25> vref<26> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X59 vref<20> vref<21> vssd sky130_fd_pr__res_generic_nd__hv w=0.29 l=350.09
X60 vddio_q vrefgen_en_h_n a_n138_3352# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X61 vssd vrefgen_en_h a_11607_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X62 a_11607_n869# vrefgen_en_h a_13320_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X63 a_13320_n869# vrefgen_en_h a_11607_n869# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
.ends

.subckt sky130_fd_io__gpiovrefv2_ctl vrefgen_en_h_n vddio_q hld_h_n enable_h selb_h<2>
+ selb_h<1> sel_h<3> sel<1> sel<3> selb_h<3> selb_h<4> sel_h<4> vrefgen_en sel<0>
+ sel<4> sel<2> sel_h<2> sel_h<1> vrefgen_en_h sel_h<0> vccd vssd selb_h<0>
Xsky130_fd_io__com_ctl_ls_0 vssd sky130_fd_io__com_ctl_ls_5/rst_h sky130_fd_io__com_ctl_ls_5/hld_h_n
+ sel<4> sel_h<4> vccd vddio_q vccd selb_h<4> vssd sky130_fd_io__com_ctl_ls
Xsky130_fd_io__com_ctl_ls_1 vssd sky130_fd_io__com_ctl_ls_5/rst_h sky130_fd_io__com_ctl_ls_5/hld_h_n
+ sel<3> sel_h<3> vccd vddio_q vccd selb_h<3> vssd sky130_fd_io__com_ctl_ls
Xsky130_fd_io__com_ctl_ls_2 vssd sky130_fd_io__com_ctl_ls_5/rst_h sky130_fd_io__com_ctl_ls_5/hld_h_n
+ sel<2> sel_h<2> vccd vddio_q vccd selb_h<2> vssd sky130_fd_io__com_ctl_ls
Xsky130_fd_io__com_ctl_ls_3 vssd sky130_fd_io__com_ctl_ls_5/rst_h sky130_fd_io__com_ctl_ls_5/hld_h_n
+ sel<1> sel_h<1> vccd vddio_q vccd selb_h<1> vssd sky130_fd_io__com_ctl_ls
Xsky130_fd_io__com_ctl_ls_4 vssd sky130_fd_io__com_ctl_ls_5/rst_h sky130_fd_io__com_ctl_ls_5/hld_h_n
+ vrefgen_en vrefgen_en_h vccd vddio_q vccd vrefgen_en_h_n vssd sky130_fd_io__com_ctl_ls
Xsky130_fd_io__com_ctl_ls_5 vssd sky130_fd_io__com_ctl_ls_5/rst_h sky130_fd_io__com_ctl_ls_5/hld_h_n
+ sel<0> sel_h<0> vccd vddio_q vccd selb_h<0> vssd sky130_fd_io__com_ctl_ls
X0 a_4618_724# hld_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X1 vssd enable_h a_5024_750# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X2 sky130_fd_io__com_ctl_ls_5/hld_h_n a_4618_724# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X3 vddio_q enable_h sky130_fd_io__com_ctl_ls_5/rst_h vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X4 a_5024_750# hld_h_n a_4618_724# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X5 sky130_fd_io__com_ctl_ls_5/hld_h_n a_4618_724# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X6 vddio_q enable_h a_4618_724# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X7 vssd enable_h sky130_fd_io__com_ctl_ls_5/rst_h vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X8 vddio_q enable_h sky130_fd_io__com_ctl_ls_5/rst_h vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X9 sky130_fd_io__com_ctl_ls_5/hld_h_n a_4618_724# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X10 a_4618_724# hld_h_n vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X11 vddio_q enable_h a_4618_724# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
.ends

.subckt sky130_fd_io__gpiovrefv2_hv_nand2 a_119_4# w_0_358# a_63_36# a_275_4# a_66_424#
+ a_219_424# VSUBS
X0 a_219_424# a_275_4# a_219_36# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0.105 ps=1.03 w=0.75 l=0.5
X1 a_219_36# a_119_4# a_63_36# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21 ps=2.06 w=0.75 l=0.5
X2 a_219_424# a_119_4# a_66_424# w_0_358# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X3 a_66_424# a_275_4# a_219_424# w_0_358# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
.ends

.subckt sky130_fd_io__gpiovrefv2_hv_inv w_0_358# a_n58_4# a_42_36# a_n114_36# a_66_424#
+ VSUBS
X0 a_42_36# a_n58_4# a_n114_36# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0.21 ps=2.06 w=0.75 l=0.5
X1 a_42_36# a_n58_4# a_66_424# w_0_358# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
.ends

.subckt sky130_fd_io__gpiovrefv2_hv_nor2 w_0_358# a_119_218# a_309_4# a_97_36# a_253_36#
+ a_219_424# VSUBS
X0 a_66_424# a_309_4# a_253_36# w_0_358# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X1 a_253_36# a_119_218# a_97_36# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21 ps=2.06 w=0.75 l=0.5
X2 a_219_424# a_119_218# a_66_424# w_0_358# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X3 a_97_36# a_309_4# a_253_36# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0.105 ps=1.03 w=0.75 l=0.5
X4 a_253_36# a_309_4# a_66_424# w_0_358# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X5 a_66_424# a_119_218# a_219_424# w_0_358# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
.ends

.subckt sky130_fd_io__gpiovrefv2_hv_nand3 a_119_4# w_0_358# a_431_4# a_63_36# a_275_4#
+ a_66_424# a_219_424# VSUBS
X0 a_219_424# a_431_4# a_375_36# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0.105 ps=1.03 w=0.75 l=0.5
X1 a_375_36# a_275_4# a_219_36# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 a_219_36# a_119_4# a_63_36# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21 ps=2.06 w=0.75 l=0.5
X3 a_219_424# a_119_4# a_66_424# w_0_358# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X4 a_219_424# a_431_4# a_66_424# w_0_358# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X5 a_66_424# a_275_4# a_219_424# w_0_358# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
.ends

.subckt sky130_fd_io__gpiovrefv2_decoder_5_32_cell vrefout vrefin vddio_q in3 in4
+ in2 in1 in0 vssd
Xsky130_fd_io__gpiovrefv2_hv_nand2_0 in4 vddio_q vssd in3 vddio_q m1_877_290# vssd
+ sky130_fd_io__gpiovrefv2_hv_nand2
Xsky130_fd_io__gpiovrefv2_hv_inv_0 vddio_q a_1853_104# a_2009_426# vssd vddio_q vssd
+ sky130_fd_io__gpiovrefv2_hv_inv
Xsky130_fd_io__gpiovrefv2_hv_nor2_0 vddio_q m1_877_290# m1_114_192# vssd a_1853_104#
+ vddio_q vssd sky130_fd_io__gpiovrefv2_hv_nor2
Xsky130_fd_io__gpiovrefv2_hv_nand3_0 in2 vddio_q in0 vssd in1 vddio_q m1_114_192#
+ vssd sky130_fd_io__gpiovrefv2_hv_nand3
X0 vrefout a_1853_104# vrefin vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1 vrefout a_1853_104# vrefin vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0.105 ps=1.03 w=0.75 l=0.5
X2 vrefout a_2009_426# vrefin vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X3 vrefin a_1853_104# vrefout vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 vrefin a_1853_104# vrefout vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21 ps=2.06 w=0.75 l=0.5
X5 vrefout a_2009_426# vrefin vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X6 vrefin a_2009_426# vrefout vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
.ends

.subckt sky130_fd_io__gpiovrefv2_decoder_5_32 vrefin vddio_q vref<30> vref<29> vref<28>
+ vref<27> vref<26> vref<25> vref<24> vref<23> vref<22> vref<21> vref<20> vref<19>
+ vref<18> vref<16> vref<15> vref<14> vref<13> vref<12> vref<11> vref<10> vref<9>
+ vref<8> vref<7> vref<6> vref<5> vref<4> vref<3> vref<2> vref<0> selb_h<4> selb_h<2>
+ selb_h<1> selb_h<0> sel_h<4> sel_h<3> sel_h<2> sel_h<1> sel_h<0> m1_0_n160# vref<1>
+ vref<17> m1_0_2532# vref<31> selb_h<3> vssd
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_1 vrefin vref<15> vddio_q sel_h<3> selb_h<4>
+ sel_h<2> sel_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_0 vrefin vref<11> vddio_q sel_h<3> selb_h<4>
+ selb_h<2> sel_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_2 vrefin vref<13> vddio_q sel_h<3> selb_h<4>
+ sel_h<2> selb_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_20 vrefin vref<20> vddio_q selb_h<3> sel_h<4>
+ sel_h<2> selb_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_31 vrefin vref<14> vddio_q sel_h<3> selb_h<4>
+ sel_h<2> sel_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_30 vrefin vref<8> vddio_q sel_h<3> selb_h<4>
+ selb_h<2> selb_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_3 vrefin vref<5> vddio_q selb_h<3> selb_h<4>
+ sel_h<2> selb_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_10 vrefin vref<29> vddio_q sel_h<3> sel_h<4>
+ sel_h<2> selb_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_21 vrefin vref<22> vddio_q selb_h<3> sel_h<4>
+ sel_h<2> sel_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_4 vrefin vref<7> vddio_q selb_h<3> selb_h<4>
+ sel_h<2> sel_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_22 vrefin vref<24> vddio_q sel_h<3> sel_h<4>
+ selb_h<2> selb_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_11 vrefin vref<19> vddio_q selb_h<3> sel_h<4>
+ selb_h<2> sel_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_5 vrefin vref<3> vddio_q selb_h<3> selb_h<4>
+ selb_h<2> sel_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_12 vrefin vref<23> vddio_q selb_h<3> sel_h<4>
+ sel_h<2> sel_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_23 vrefin vref<16> vddio_q selb_h<3> sel_h<4>
+ selb_h<2> selb_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_6 vrefin vref<1> vddio_q selb_h<3> selb_h<4>
+ selb_h<2> selb_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_13 vrefin vref<21> vddio_q selb_h<3> sel_h<4>
+ sel_h<2> selb_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_7 vrefin vref<9> vddio_q sel_h<3> selb_h<4>
+ selb_h<2> selb_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_24 vrefin vref<4> vddio_q selb_h<3> selb_h<4>
+ sel_h<2> selb_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_14 vrefin vref<31> vddio_q sel_h<3> sel_h<4>
+ sel_h<2> sel_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_8 vrefin vref<25> vddio_q sel_h<3> sel_h<4>
+ selb_h<2> selb_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_25 vrefin vref<0> vddio_q selb_h<3> selb_h<4>
+ selb_h<2> selb_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_9 vrefin vref<27> vddio_q sel_h<3> sel_h<4>
+ selb_h<2> sel_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_15 vrefin vref<17> vddio_q selb_h<3> sel_h<4>
+ selb_h<2> selb_h<1> sel_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_26 vrefin vref<6> vddio_q selb_h<3> selb_h<4>
+ sel_h<2> sel_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_16 vrefin vref<30> vddio_q sel_h<3> sel_h<4>
+ sel_h<2> sel_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_27 vrefin vref<2> vddio_q selb_h<3> selb_h<4>
+ selb_h<2> sel_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_18 vrefin vref<26> vddio_q sel_h<3> sel_h<4>
+ selb_h<2> sel_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_17 vrefin vref<18> vddio_q selb_h<3> sel_h<4>
+ selb_h<2> sel_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_28 vrefin vref<12> vddio_q sel_h<3> selb_h<4>
+ sel_h<2> selb_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_29 vrefin vref<10> vddio_q sel_h<3> selb_h<4>
+ selb_h<2> sel_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
Xsky130_fd_io__gpiovrefv2_decoder_5_32_cell_19 vrefin vref<28> vddio_q sel_h<3> sel_h<4>
+ sel_h<2> selb_h<1> selb_h<0> vssd sky130_fd_io__gpiovrefv2_decoder_5_32_cell
.ends

.subckt sky130_fd_io__top_gpiovrefv2 ref_sel<4> ref_sel<3> ref_sel<1> vrefgen_en hld_h_n
+ enable_h ref_sel<2> ref_sel<0> vinref vddio_q vddio vssio vssa vccd vcchib vswitch
+ vssio_q vdda vssd amuxbus_b amuxbus_a
Xsky130_fd_io__gpiovrefv2_res_ladder_0 sky130_fd_io__gpiovrefv2_ctl_0/vrefgen_en_h
+ sky130_fd_io__gpiovrefv2_ctl_0/vrefgen_en_h_n sky130_fd_io__gpiovrefv2_res_ladder_0/vref<31>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<30> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<29>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<28> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<27>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<26> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<25>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<24> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<23>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<22> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<21>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<20> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<19>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<18> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<17>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<16> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<15>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<14> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<13>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<12> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<11>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<10> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<9>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<8> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<7>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<6> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<5>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<4> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<3>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<2> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<1>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<0> vssd vddio_q vssd vssd sky130_fd_io__gpiovrefv2_res_ladder
Xsky130_fd_io__gpiovrefv2_ctl_0 sky130_fd_io__gpiovrefv2_ctl_0/vrefgen_en_h_n vddio_q
+ hld_h_n enable_h sky130_fd_io__gpiovrefv2_ctl_0/selb_h<2> sky130_fd_io__gpiovrefv2_ctl_0/selb_h<1>
+ sky130_fd_io__gpiovrefv2_ctl_0/sel_h<3> ref_sel<1> ref_sel<3> sky130_fd_io__gpiovrefv2_ctl_0/selb_h<3>
+ sky130_fd_io__gpiovrefv2_ctl_0/selb_h<4> sky130_fd_io__gpiovrefv2_ctl_0/sel_h<4>
+ vrefgen_en ref_sel<0> ref_sel<4> ref_sel<2> sky130_fd_io__gpiovrefv2_ctl_0/sel_h<2>
+ sky130_fd_io__gpiovrefv2_ctl_0/sel_h<1> sky130_fd_io__gpiovrefv2_ctl_0/vrefgen_en_h
+ sky130_fd_io__gpiovrefv2_ctl_0/sel_h<0> vccd vssd sky130_fd_io__gpiovrefv2_ctl_0/selb_h<0>
+ sky130_fd_io__gpiovrefv2_ctl
Xsky130_fd_io__gpiovrefv2_decoder_5_32_0 vinref vddio_q sky130_fd_io__gpiovrefv2_res_ladder_0/vref<30>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<29> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<28>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<27> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<26>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<25> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<24>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<23> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<22>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<21> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<20>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<19> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<18>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<16> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<15>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<14> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<13>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<12> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<11>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<10> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<9>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<8> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<7>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<6> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<5>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<4> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<3>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<2> sky130_fd_io__gpiovrefv2_res_ladder_0/vref<0>
+ sky130_fd_io__gpiovrefv2_ctl_0/selb_h<4> sky130_fd_io__gpiovrefv2_ctl_0/selb_h<2>
+ sky130_fd_io__gpiovrefv2_ctl_0/selb_h<1> sky130_fd_io__gpiovrefv2_ctl_0/selb_h<0>
+ sky130_fd_io__gpiovrefv2_ctl_0/sel_h<4> sky130_fd_io__gpiovrefv2_ctl_0/sel_h<3>
+ sky130_fd_io__gpiovrefv2_ctl_0/sel_h<2> sky130_fd_io__gpiovrefv2_ctl_0/sel_h<1>
+ sky130_fd_io__gpiovrefv2_ctl_0/sel_h<0> vssd sky130_fd_io__gpiovrefv2_res_ladder_0/vref<1>
+ sky130_fd_io__gpiovrefv2_res_ladder_0/vref<17> vssd sky130_fd_io__gpiovrefv2_res_ladder_0/vref<31>
+ sky130_fd_io__gpiovrefv2_ctl_0/selb_h<3> vssd sky130_fd_io__gpiovrefv2_decoder_5_32
X0 vssd sky130_fd_io__gpiovrefv2_ctl_0/vrefgen_en_h_n vinref vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X1 vinref sky130_fd_io__gpiovrefv2_ctl_0/vrefgen_en_h_n vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
.ends

.subckt sky130_ef_io__vssa_hvc_clamped_pad VSSD VSSA VDDIO VSSA_PAD VSWITCH VSSIO
+ VCCHIB VDDA VDDIO_Q AMUXBUS_A AMUXBUS_B VSSIO_Q VCCD
Xsky130_fd_io__top_ground_hvc_wpad_0 VCCHIB VDDA VDDIO_Q VSSIO_Q VSSA_PAD sky130_fd_io__top_ground_hvc_wpad_0/PADISOR
+ sky130_fd_io__top_ground_hvc_wpad_0/PADISOL VDDA VSSA VDDIO VSSA AMUXBUS_B VSSIO
+ VDDIO VSSD VSWITCH VSSA AMUXBUS_A VCCD sky130_fd_io__top_ground_hvc_wpad
.ends

.subckt chip_io_gpio_connects_vert tie_lo_esd pad_a_esd_1_h dm[1] dm[0] analog_pol
+ inp_dis enable_h hld_h_n dm[2] hld_ovr out enable_vswitch_h enable_vdda_h vtrip_sel
+ oe_n tie_hi_esd in enable_vddio slow pad_a_esd_0_h pad_a_noesd_h analog_en analog_sel
+ ib_mode_sel in_h zero one enable_inp_h constant_block_0/vccd VSUBS
Xconstant_block_0 one constant_block_0/vccd zero VSUBS constant_block
.ends

.subckt s8_esd_res75only_small pad rout
X0 pad rout sky130_fd_pr__res_generic_po w=2 l=3.15
.ends

.subckt sky130_fd_io__amuxsplitv2_switch pgate_sl_h_n pgate_sr_h_n ngate_sl_h ngate_sr_h
+ nmid_h amuxbus_l amuxbus_r vdda vssa w_4833_342#
Xs8_esd_res75only_small_0 vssa s8_esd_res75only_small_0/rout s8_esd_res75only_small
X0 w_4833_342# pgate_sl_h_n amuxbus_l vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X1 amuxbus_r pgate_sr_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X2 amuxbus_l pgate_sl_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X3 amuxbus_r pgate_sr_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X4 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X5 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X6 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X7 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X8 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X9 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X10 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X11 amuxbus_l pgate_sl_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X12 w_4833_342# pgate_sr_h_n amuxbus_r vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X13 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X14 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X15 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X16 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X17 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X18 w_4833_342# pgate_sr_h_n amuxbus_r vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X19 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X20 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X21 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X22 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X23 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X24 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X25 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=2.8 ps=20.56 w=10 l=0.5
X26 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X27 w_4833_342# pgate_sr_h_n amuxbus_r vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X28 amuxbus_r pgate_sr_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X29 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X30 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X31 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X32 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X33 w_4833_342# pgate_sl_h_n amuxbus_l vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X34 amuxbus_l pgate_sl_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X35 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X36 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X37 w_4833_342# pgate_sr_h_n amuxbus_r vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X38 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X39 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X40 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X41 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X42 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X43 w_4833_342# pgate_sl_h_n amuxbus_l vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X44 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X45 amuxbus_r pgate_sr_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X46 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=2.8 ps=20.56 w=10 l=0.5
X47 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X48 w_4833_342# pgate_sr_h_n amuxbus_r vdda sky130_fd_pr__pfet_g5v0d10v5 ad=2.8 pd=20.56 as=1.4 ps=10.28 w=10 l=0.5
X49 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X50 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=2.8 pd=20.56 as=1.4 ps=10.28 w=10 l=0.5
X51 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X52 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X53 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X54 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X55 amuxbus_l pgate_sl_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X56 w_4833_342# pgate_sl_h_n amuxbus_l vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X57 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X58 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X59 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X60 amuxbus_r pgate_sr_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X61 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X62 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X63 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X64 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X65 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X66 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X67 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X68 amuxbus_l pgate_sl_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=2.8 ps=20.56 w=10 l=0.5
X69 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X70 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X71 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X72 w_4833_342# pgate_sl_h_n amuxbus_l vdda sky130_fd_pr__pfet_g5v0d10v5 ad=2.8 pd=20.56 as=1.4 ps=10.28 w=10 l=0.5
X73 w_4833_342# pgate_sl_h_n amuxbus_l vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X74 amuxbus_l pgate_sl_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X75 amuxbus_l pgate_sl_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X76 amuxbus_r pgate_sr_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=2.8 ps=20.56 w=10 l=0.5
X77 w_4833_342# pgate_sr_h_n amuxbus_r vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X78 w_4833_342# nmid_h s8_esd_res75only_small_0/rout vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.56 w=5 l=0.5
X79 amuxbus_l ngate_sl_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X80 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X81 amuxbus_r pgate_sr_h_n w_4833_342# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X82 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X83 w_4833_342# pgate_sl_h_n amuxbus_l vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X84 s8_esd_res75only_small_0/rout nmid_h w_4833_342# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.56 as=0.7 ps=5.28 w=5 l=0.5
X85 w_4833_342# ngate_sl_h amuxbus_l w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X86 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=2.8 pd=20.56 as=1.4 ps=10.28 w=10 l=0.5
X87 w_4833_342# ngate_sr_h amuxbus_r w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X88 w_4833_342# pgate_sr_h_n amuxbus_r vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
X89 amuxbus_r ngate_sr_h w_4833_342# w_4833_342# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.28 as=1.4 ps=10.28 w=10 l=0.5
.ends

.subckt sky130_fd_io__top_amuxsplitv2 amuxbus_a_r amuxbus_a_l amuxbus_b_r amuxbus_b_l
+ enable_vdda_h hld_vdda_h_n switch_aa_s0 switch_aa_sl switch_aa_sr switch_bb_s0 switch_bb_sl
+ switch_bb_sr vssd vssio vswitch vccd vddio_q vddio vcchib w_2174_29699# w_2174_23399#
+ vdda vssa vssio_q
Xsky130_fd_io__amuxsplitv2_switch_1 sky130_fd_io__amuxsplitv2_switch_1/pgate_sl_h_n
+ sky130_fd_io__amuxsplitv2_switch_1/pgate_sr_h_n sky130_fd_io__amuxsplitv2_switch_1/ngate_sl_h
+ sky130_fd_io__amuxsplitv2_switch_1/ngate_sr_h sky130_fd_io__amuxsplitv2_switch_1/nmid_h
+ amuxbus_a_l amuxbus_a_r vdda vssa w_2174_29699# sky130_fd_io__amuxsplitv2_switch
Xsky130_fd_io__amuxsplitv2_switch_0 sky130_fd_io__amuxsplitv2_switch_0/pgate_sl_h_n
+ sky130_fd_io__amuxsplitv2_switch_0/pgate_sr_h_n sky130_fd_io__amuxsplitv2_switch_0/ngate_sl_h
+ sky130_fd_io__amuxsplitv2_switch_0/ngate_sr_h sky130_fd_io__amuxsplitv2_switch_0/nmid_h
+ amuxbus_b_l amuxbus_b_r vdda vssa w_2174_23399# sky130_fd_io__amuxsplitv2_switch
X0 a_6162_10251# vccd a_5456_10673# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 a_6492_10251# vccd a_5456_10959# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X2 vssa a_5554_2103# a_5498_2867# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X3 a_3092_13912# a_3060_13812# vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X4 vssa a_2990_15060# a_6492_14039# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 vssa a_3060_13144# sky130_fd_io__amuxsplitv2_switch_0/ngate_sl_h vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X6 a_3060_8764# a_5358_3495# a_5456_8758# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X7 a_5554_2103# a_6187_2069# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X8 vssa a_2990_4191# a_6492_3675# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 vssa a_2990_4964# a_6492_5203# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10 sky130_fd_io__amuxsplitv2_switch_1/pgate_sl_h_n a_3060_6506# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X11 a_3092_8864# a_5358_3495# a_5456_9044# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X12 a_3060_8096# a_3092_8329# vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X13 a_3092_13377# a_5325_2867# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 vssa a_2958_11981# a_6162_12775# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 sky130_fd_io__amuxsplitv2_switch_0/pgate_sl_h_n a_3060_11554# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X16 a_5456_9044# vccd a_6162_8991# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X17 vdda a_3060_15668# sky130_fd_io__amuxsplitv2_switch_0/pgate_sr_h_n vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X18 vssa a_2990_15060# a_6492_14039# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_6162_10251# vccd a_5456_10673# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X20 a_6492_10251# vccd a_5456_10959# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X21 a_6492_8991# a_2990_10012# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X22 a_6768_2037# hld_vdda_h_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X23 a_6492_5203# vccd a_5456_5911# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X24 a_6162_15299# vccd a_5456_15721# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X25 a_6492_15299# vccd a_5456_16007# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X26 vssa a_2958_11981# a_6162_12775# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 vdda a_3060_15954# a_3060_15668# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X28 vssa a_2958_11981# a_6162_11515# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X29 a_3092_5805# a_5325_2867# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X30 a_6162_7727# a_2958_6933# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X31 vssa a_2958_11981# a_6162_11515# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 vssa a_2990_10012# a_6492_10251# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X33 vswitch a_3092_8864# a_3060_8764# vswitch sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X34 vdda a_5554_2103# a_5325_2867# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X35 a_5456_6520# vccd a_6162_6467# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X36 vssa a_2990_12031# a_6492_11515# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X37 vssa a_2990_10012# a_6492_10251# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X38 a_6162_6467# a_2958_6933# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X39 a_6492_12775# vccd a_5456_13483# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X40 vssa a_3060_10620# sky130_fd_io__amuxsplitv2_switch_1/pgate_sr_h_n vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X41 a_6492_3675# vccd a_5456_3442# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X42 a_6162_12775# vccd a_5456_13197# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X43 vssa a_2958_9962# a_6162_10251# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X44 a_6162_6467# a_2958_6933# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X45 a_2990_12031# a_2958_11981# vssd vssd sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X46 vdda enable_vdda_h a_6187_2069# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X47 vssd switch_bb_sr a_2958_15010# vssd sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X48 vssd switch_bb_s0 a_2958_4914# vssd sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X49 vccd a_2958_4141# a_2990_4191# vccd sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X50 a_6162_14039# vccd a_5456_14092# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X51 a_6492_14039# vccd a_5456_13806# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X52 a_6492_8991# vccd a_5456_8758# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X53 a_6492_5203# a_2990_4964# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X54 vccd switch_aa_sr a_2958_9962# vccd sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X55 a_6162_5203# a_2958_4914# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X56 vdda a_3092_3548# a_3060_3448# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X57 a_5554_2103# a_6187_2069# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X58 a_6492_3675# vccd a_5456_3442# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X59 a_5456_6234# vccd a_6492_6467# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X60 vssa a_3060_15668# sky130_fd_io__amuxsplitv2_switch_0/pgate_sr_h_n vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X61 vssa a_5325_2867# a_3060_6506# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X62 vssa a_5325_2867# a_3092_13912# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X63 a_5358_3495# a_5325_2867# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X64 a_2990_4964# a_2958_4914# vccd vccd sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X65 a_5456_10959# a_5358_3495# a_3060_10906# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X66 a_2958_4141# switch_aa_s0 vssd vssd sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X67 a_3060_15668# a_5325_2867# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X68 a_3060_10906# a_3060_10620# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X69 a_6492_11515# a_2990_12031# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X70 a_6162_12775# vccd a_5456_13197# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X71 a_6492_12775# vccd a_5456_13483# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X72 a_5456_5625# vccd a_6162_5203# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X73 a_6492_11515# a_2990_12031# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X74 vssa a_2958_4141# a_6162_3675# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X75 a_6162_6467# vccd a_5456_6520# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X76 a_5456_10673# vccd a_6162_10251# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X77 a_5456_10959# vccd a_6492_10251# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X78 a_5456_5911# vccd a_6492_5203# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X79 a_6162_10251# a_2958_9962# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X80 sky130_fd_io__amuxsplitv2_switch_1/pgate_sl_h_n a_3060_6506# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X81 vssa a_2958_15010# a_6162_14039# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X82 vdda a_3060_5572# a_3092_5805# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X83 a_6492_8991# a_2990_10012# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X84 a_5364_2361# a_6768_2037# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X85 a_2958_11981# switch_bb_sl vssd vssd sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X86 a_6162_8991# a_2958_9962# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X87 vssa enable_vdda_h a_6187_2069# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X88 a_6162_6467# vccd a_5456_6520# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X89 a_6162_7727# a_2958_6933# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X90 a_6162_8991# a_2958_9962# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X91 a_5456_3728# vccd a_6162_3675# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X92 a_5456_8149# vccd a_6162_7727# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X93 a_6492_7727# a_2990_6983# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X94 a_2990_6983# a_2958_6933# vssd vssd sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X95 a_3060_3448# a_5358_3495# a_5456_3442# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X96 a_6162_3675# a_2958_4141# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X97 a_6492_7727# a_2990_6983# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X98 vssa a_3060_5572# sky130_fd_io__amuxsplitv2_switch_0/nmid_h vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X99 a_3060_11288# a_5358_3495# a_5456_11282# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X100 a_5456_8758# vccd a_6492_8991# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X101 a_6492_3675# a_2990_4191# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X102 a_3092_3548# a_5358_3495# a_5456_3728# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X103 a_6492_15299# a_2990_15060# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X104 a_6492_14039# a_2990_15060# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X105 a_5358_3495# a_5325_2867# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X106 a_6492_3675# a_2990_4191# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X107 a_6492_5203# a_2990_4964# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X108 a_3060_11554# a_5358_3495# a_5456_11568# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X109 a_6162_5203# vccd a_5456_5625# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X110 sky130_fd_io__amuxsplitv2_switch_1/ngate_sr_h a_3060_8764# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X111 vdda a_6187_2069# a_5554_2103# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X112 a_5456_8758# vccd a_6492_8991# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X113 vdda a_6768_2037# a_5364_2361# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X114 a_5456_3728# vccd a_6162_3675# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X115 a_5456_11568# vccd a_6162_11515# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X116 a_5456_11282# vccd a_6492_11515# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X117 a_5456_8149# vccd a_6162_7727# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X118 a_6162_8991# vccd a_5456_9044# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X119 a_2990_15060# a_2958_15010# vccd vccd sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X120 a_5364_2361# a_6768_2037# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X121 sky130_fd_io__amuxsplitv2_switch_0/pgate_sl_h_n a_3060_11554# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X122 a_6162_11515# a_2958_11981# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X123 vccd a_2958_11981# a_2990_12031# vccd sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X124 vdda a_3060_10906# a_3060_10620# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X125 vssa a_2958_6933# a_6162_6467# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X126 a_5456_6234# vccd a_6492_6467# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X127 vssa a_2990_15060# a_6492_15299# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X128 vssa a_3060_8096# sky130_fd_io__amuxsplitv2_switch_1/ngate_sl_h vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X129 a_2958_4141# switch_aa_s0 vccd vccd sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X130 a_3060_13812# a_5358_3495# a_5456_13806# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X131 a_5456_10673# a_5358_3495# a_3060_10620# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X132 a_6162_10251# a_2958_9962# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X133 vssa a_2990_6983# a_6492_6467# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X134 vssa a_2958_15010# a_6162_15299# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X135 vssa a_2990_4964# a_6492_5203# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X136 sky130_fd_io__amuxsplitv2_switch_1/ngate_sr_h a_3060_8764# vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X137 vssa a_2990_6983# a_6492_6467# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X138 a_3092_8329# a_5325_2867# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X139 vssa a_2958_15010# a_6162_15299# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X140 vssa a_2958_4914# a_6162_5203# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X141 a_6162_7727# vccd a_5456_8149# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X142 a_5456_11568# vccd a_6162_11515# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X143 a_5456_11282# vccd a_6492_11515# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X144 sky130_fd_io__amuxsplitv2_switch_1/nmid_h a_3060_3448# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X145 vssa a_2958_4914# a_6162_5203# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X146 vdda a_3060_5572# sky130_fd_io__amuxsplitv2_switch_0/nmid_h vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X147 vccd switch_bb_s0 a_2958_4914# vccd sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X148 vssa a_2958_15010# a_6162_14039# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X149 a_5456_10673# vccd a_6162_10251# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X150 a_5456_10959# vccd a_6492_10251# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X151 a_3060_5572# a_3092_5805# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X152 a_3092_13912# a_5358_3495# a_5456_14092# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X153 vssa a_6187_2069# a_5554_2103# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X154 vdda a_3060_11554# a_3060_11288# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X155 vssa a_2990_12031# a_6492_12775# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X156 vssa a_6768_2037# a_5364_2361# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X157 vccd switch_bb_sr a_2958_15010# vccd sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X158 vssa a_2990_12031# a_6492_12775# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X159 a_5456_14092# vccd a_6162_14039# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X160 a_5456_13806# vccd a_6492_14039# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X161 a_5456_5911# vccd a_6492_5203# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X162 a_2958_11981# switch_bb_sl vccd vccd sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X163 a_6492_11515# vccd a_5456_11282# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X164 a_6162_7727# vccd a_5456_8149# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X165 vssd a_2958_9962# a_2990_10012# vssd sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X166 a_6162_11515# vccd a_5456_11568# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X167 a_6492_6467# vccd a_5456_6234# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X168 sky130_fd_io__amuxsplitv2_switch_0/ngate_sr_h a_3060_13812# vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X169 vssa a_2990_10012# a_6492_8991# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X170 vccd a_2958_6933# a_2990_6983# vccd sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X171 a_5456_14092# vccd a_6162_14039# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X172 a_5456_13806# vccd a_6492_14039# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X173 a_2958_6933# switch_aa_sl vssd vssd sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X174 a_6162_15299# vccd a_5456_15721# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X175 a_6492_15299# vccd a_5456_16007# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X176 vssa a_2958_6933# a_6162_7727# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X177 a_5456_13197# a_5358_3495# a_3092_13377# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X178 vssa a_5325_2867# a_3092_8864# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X179 vssa a_2990_10012# a_6492_8991# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X180 a_6162_3675# a_2958_4141# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X181 a_6162_11515# vccd a_5456_11568# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X182 a_6492_11515# vccd a_5456_11282# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X183 a_5456_3442# vccd a_6492_3675# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X184 a_6162_5203# vccd a_5456_5625# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X185 a_6492_6467# vccd a_5456_6234# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X186 a_3060_6506# a_3060_6240# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X187 a_6162_14039# a_2958_15010# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X188 a_5456_13197# vccd a_6162_12775# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X189 a_5456_13483# vccd a_6492_12775# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X190 a_5456_8435# vccd a_6492_7727# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X191 a_5456_13483# a_5358_3495# a_3060_13144# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X192 a_6162_12775# a_2958_11981# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X193 vssa a_5325_2867# a_3092_3548# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X194 vssa a_2958_6933# a_6162_6467# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X195 a_3060_13144# a_3092_13377# vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X196 vssa a_2990_15060# a_6492_15299# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X197 a_6492_14039# a_2990_15060# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X198 a_5456_5625# a_5358_3495# a_3092_5805# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X199 a_6162_12775# a_2958_11981# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X200 vswitch a_3060_8096# sky130_fd_io__amuxsplitv2_switch_1/ngate_sl_h vswitch sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X201 a_6162_11515# a_2958_11981# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X202 vdda a_3060_10620# sky130_fd_io__amuxsplitv2_switch_1/pgate_sr_h_n vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X203 a_6162_14039# vccd a_5456_14092# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X204 a_6492_14039# vccd a_5456_13806# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X205 a_6162_3675# vccd a_5456_3728# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X206 vswitch a_3060_8096# a_3092_8329# vswitch sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X207 a_6492_10251# a_2990_10012# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X208 a_6492_5203# vccd a_5456_5911# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X209 vswitch a_3092_13912# a_3060_13812# vswitch sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X210 a_6492_10251# a_2990_10012# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X211 sky130_fd_io__amuxsplitv2_switch_1/nmid_h a_3060_3448# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X212 vssd switch_aa_sr a_2958_9962# vssd sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X213 a_6162_8991# vccd a_5456_9044# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X214 a_5456_13483# vccd a_6492_12775# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X215 a_5456_8435# vccd a_6492_7727# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X216 a_5456_3442# vccd a_6492_3675# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X217 a_5456_13197# vccd a_6162_12775# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X218 a_6162_3675# vccd a_5456_3728# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X219 a_5456_6520# vccd a_6162_6467# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X220 vssd a_2958_4914# a_2990_4964# vssd sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X221 a_6492_8991# vccd a_5456_8758# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X222 a_5325_2867# a_5364_2361# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X223 a_3060_11554# a_3060_11288# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X224 a_2990_10012# a_2958_9962# vccd vccd sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X225 a_3092_8864# a_3060_8764# vswitch vswitch sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X226 a_5456_16007# a_5358_3495# a_3060_15954# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X227 a_3060_6240# a_5358_3495# a_5456_6234# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X228 a_3060_15954# a_3060_15668# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X229 a_6492_15299# a_2990_15060# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X230 a_3060_10620# a_5325_2867# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X231 a_6492_6467# a_2990_6983# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X232 a_3060_6506# a_5358_3495# a_5456_6520# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X233 a_5456_15721# a_5358_3495# a_3060_15668# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X234 a_6162_15299# a_2958_15010# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X235 a_5456_15721# vccd a_6162_15299# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X236 a_5456_16007# vccd a_6492_15299# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X237 a_5498_2867# a_5364_2361# a_5325_2867# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X238 a_6492_6467# a_2990_6983# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X239 a_6162_15299# a_2958_15010# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X240 a_2990_4191# a_2958_4141# vssd vssd sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X241 a_5456_5625# vccd a_6162_5203# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X242 vssa a_2990_12031# a_6492_11515# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X243 a_6768_2037# hld_vdda_h_n vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X244 a_6162_5203# a_2958_4914# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X245 a_6492_7727# vccd a_5456_8435# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X246 a_3092_3548# a_3060_3448# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X247 a_5456_8149# a_5358_3495# a_3092_8329# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X248 vssa a_2958_9962# a_6162_10251# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X249 a_6162_14039# a_2958_15010# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X250 vswitch a_3060_13144# sky130_fd_io__amuxsplitv2_switch_0/ngate_sl_h vswitch sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X251 a_5456_15721# vccd a_6162_15299# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X252 a_5456_16007# vccd a_6492_15299# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X253 a_5456_8435# a_5358_3495# a_3060_8096# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X254 sky130_fd_io__amuxsplitv2_switch_0/ngate_sr_h a_3060_13812# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X255 a_6492_12775# a_2990_12031# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X256 vssa a_2958_9962# a_6162_8991# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X257 vswitch a_3060_13144# a_3092_13377# vswitch sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X258 vdda a_5554_2103# a_5325_2867# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X259 a_6492_12775# a_2990_12031# vssa vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X260 vssa a_2958_9962# a_6162_8991# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X261 vssa a_2990_6983# a_6492_7727# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X262 a_5325_2867# a_5364_2361# vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X263 vdda a_3060_6506# a_3060_6240# vdda sky130_fd_pr__pfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X264 vssa a_5325_2867# a_3060_11554# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X265 vssa a_2958_4141# a_6162_3675# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X266 a_5456_5911# a_5358_3495# a_3060_5572# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X267 vssa a_2990_6983# a_6492_7727# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X268 a_5456_9044# vccd a_6162_8991# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X269 vssd a_2958_15010# a_2990_15060# vssd sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X270 a_2958_6933# switch_aa_sl vccd vccd sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
X271 vssa a_2990_4191# a_6492_3675# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X272 vssa a_2958_6933# a_6162_7727# vssa sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X273 a_6492_7727# vccd a_5456_8435# vssa sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
.ends

.subckt sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad vcc_io a_10282_1285# a_5322_1285#
+ a_8980_1457# a_7988_1457# a_2036_1457# a_13940_1457# a_12948_1457# a_12266_1285#
+ a_7306_1285# a_5012_1457# a_3900_1285# a_2908_1285# a_5884_1285# a_14178_1285# a_10844_1285#
+ a_1354_1285# a_7868_1285# a_12828_1285# a_8860_1285# a_13820_1285# a_4330_1285#
+ a_3338_1285# a_6996_1457# a_11956_1457# a_1044_1457# a_11274_1285# a_6314_1285#
+ a_9972_1457# a_4020_1457# a_3028_1457# a_8298_1285# w_362_785# a_13258_1285# a_9290_1285#
+ a_1916_1285# a_6004_1457# a_4892_1285# a_6876_1285# a_924_1285# a_11836_1285# a_2346_1285#
+ a_9852_1285# a_10964_1457#
X0 a_10964_1457# a_10844_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X1 a_9972_1457# a_9852_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X2 w_362_785# a_2346_1285# a_2036_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X3 a_2036_1457# a_1916_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X4 a_6996_1457# a_6876_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X5 w_362_785# a_12266_1285# a_11956_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X6 w_362_785# a_6314_1285# a_6004_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X7 a_11956_1457# a_11836_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X8 w_362_785# a_9290_1285# a_8980_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X9 a_5012_1457# a_4892_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X10 w_362_785# a_4330_1285# a_4020_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X11 a_8980_1457# a_8860_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X12 w_362_785# a_10282_1285# a_9972_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X13 w_362_785# a_3338_1285# a_3028_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X14 w_362_785# a_8298_1285# a_7988_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X15 a_1044_1457# a_924_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.425 ps=11.37 w=5 l=0.6
X16 a_4020_1457# a_3900_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X17 a_13940_1457# a_13820_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=2.975 pd=6.19 as=3.775 ps=11.51 w=5 l=0.6
X18 a_3028_1457# a_2908_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X19 a_7988_1457# a_7868_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X20 w_362_785# a_13258_1285# a_12948_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X21 w_362_785# a_7306_1285# a_6996_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X22 a_12948_1457# a_12828_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X23 w_362_785# a_14178_1285# a_13940_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.425 pd=11.37 as=2.975 ps=6.19 w=5 l=0.6
X24 w_362_785# a_1354_1285# a_1044_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X25 a_6004_1457# a_5884_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X26 w_362_785# a_11274_1285# a_10964_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X27 w_362_785# a_5322_1285# a_5012_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X28 a_9972_1457# a_9852_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X29 a_10964_1457# a_10844_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X30 w_362_785# a_2346_1285# a_2036_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X31 a_6996_1457# a_6876_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X32 w_362_785# a_6314_1285# a_6004_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X33 a_2036_1457# a_1916_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X34 w_362_785# a_12266_1285# a_11956_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X35 a_11956_1457# a_11836_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X36 a_5012_1457# a_4892_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X37 w_362_785# a_9290_1285# a_8980_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X38 a_8980_1457# a_8860_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X39 w_362_785# a_10282_1285# a_9972_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X40 w_362_785# a_4330_1285# a_4020_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X41 a_1044_1457# a_924_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.425 ps=11.37 w=5 l=0.6
X42 a_4020_1457# a_3900_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X43 w_362_785# a_3338_1285# a_3028_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X44 w_362_785# a_8298_1285# a_7988_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X45 a_3028_1457# a_2908_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X46 a_7988_1457# a_7868_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X47 w_362_785# a_7306_1285# a_6996_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X48 a_13940_1457# a_13820_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=2.975 pd=6.19 as=3.775 ps=11.51 w=5 l=0.6
X49 w_362_785# a_13258_1285# a_12948_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X50 a_12948_1457# a_12828_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X51 w_362_785# a_1354_1285# a_1044_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X52 w_362_785# a_14178_1285# a_13940_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.425 pd=11.37 as=2.975 ps=6.19 w=5 l=0.6
X53 a_6004_1457# a_5884_1285# w_362_785# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X54 w_362_785# a_5322_1285# a_5012_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X55 w_362_785# a_11274_1285# a_10964_1457# w_362_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
.ends

.subckt sky130_fd_io__top_analog_pad_pddrvr_strong vgnd_io tie_lo_esd force_lo_h pd_h<3>
+ pd_h<2> force_lovol_h vssio_amx vcc_io sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_2036_1457#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_12948_1457# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_13940_1457#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_5012_1457# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_6996_1457#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_1044_1457# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_11956_1457#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_9972_1457# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_3028_1457#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_4020_1457# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_6004_1457#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_10964_1457# w_290_3254# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_7988_1457#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_8980_1457#
Xsky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0 vcc_io pd_h<3> m1_9769_3898#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_8980_1457# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_7988_1457#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_2036_1457# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_13940_1457#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_12948_1457# m1_2697_3898#
+ m1_7657_3898# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_5012_1457# m1_11193_3898#
+ m1_11193_3898# m1_8232_3898# m1_785_3898# pd_h<3> m1_12747_3898# pd_h<2> m1_2135_3898#
+ pd_h<2> m1_785_3898# m1_9769_3898# m1_11193_3898# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_6996_1457#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_11956_1457# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_1044_1457#
+ pd_h<3> m1_8232_3898# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_9972_1457#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_4020_1457# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_3028_1457#
+ pd_h<2> w_290_3254# m1_785_3898# pd_h<3> m1_12747_3898# sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_6004_1457#
+ m1_9769_3898# m1_8232_3898# m1_12747_3898# pd_h<3> m1_12747_3898# pd_h<3> sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad_0/a_10964_1457#
+ sky130_fd_io__NFET_con_diff_wo_abt_270_analog_pad
R0 m2_413_900# tie_lo_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R1 m2_7664_899# tie_lo_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 m2_10415_900# pd_h<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R3 m2_9366_899# tie_lo_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 m1_2697_3898# m2_2790_900# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 m2_2790_900# pd_h<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R6 m2_11329_899# pd_h<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 m1_2135_3898# m2_1848_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 m2_10846_899# tie_lo_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 m1_7657_3898# m2_6804_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 m1_12747_3898# m2_12763_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 m1_12747_3898# m2_13622_900# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 m2_11758_900# pd_h<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 m1_2135_3898# m2_1260_900# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 m2_1260_900# pd_h<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 m1_785_3898# m2_897_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X0 tie_lo_esd vgnd_io sky130_fd_pr__res_generic_po w=0.5 l=10.2
R16 m2_12763_899# pd_h<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 m2_6804_899# pd_h<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R18 m1_11193_3898# m2_12189_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 m2_8506_899# pd_h<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m1_9769_3898# m2_9986_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 m1_785_3898# m2_413_900# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 m1_2697_3898# m2_3095_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R23 m1_8232_3898# m2_9366_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 m2_1565_899# pd_h<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 m2_8935_900# pd_h<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 m2_1848_899# tie_lo_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 m2_3095_899# pd_h<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 m1_11193_3898# m2_11758_900# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R29 m2_12189_899# tie_lo_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R30 m1_8232_3898# m2_8935_900# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R31 m1_9769_3898# m2_10846_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R32 m2_13622_900# tie_lo_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R33 m1_785_3898# m2_656_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R34 m1_11193_3898# m2_11329_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R35 m2_656_899# pd_h<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R36 m2_3378_899# tie_lo_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R37 m1_2135_3898# m2_1565_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R38 m1_2697_3898# m2_3378_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R39 m1_8232_3898# m2_8506_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R40 m1_9769_3898# m2_10415_900# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R41 m2_897_899# pd_h<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R42 m2_13193_899# pd_h<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R43 m1_7657_3898# m2_7664_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R44 m2_7233_900# pd_h<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R45 m1_7657_3898# m2_7233_900# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R46 m1_12747_3898# m2_13193_1200# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R47 m2_9986_899# pd_h<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad w_415_600# a_4969_1552#
+ a_2303_1380# a_5961_1552# a_13777_1380# a_8817_1380# a_4287_1380# a_10921_1552#
+ a_7945_1552# a_12905_1552# a_7263_1380# a_12223_1380# a_9929_1552# a_9247_1380#
+ a_2865_1380# a_1993_1552# a_5841_1380# a_4849_1380# a_10801_1380# a_14135_1380#
+ a_1311_1380# a_3977_1552# a_12785_1380# a_7825_1380# a_3295_1380# a_6953_1552# a_9809_1380#
+ a_11913_1552# a_1001_1552# a_6271_1380# a_5279_1380# a_11231_1380# a_10239_1380#
+ a_13897_1552# a_8937_1552# a_8255_1380# a_1873_1380# a_13215_1380# a_3857_1380#
+ a_2985_1552# a_11793_1380# a_881_1380# a_6833_1380#
X0 a_13897_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.975 pd=6.19 as=3.775 ps=11.51 w=5 l=0.6
X1 w_415_600# a_10239_1380# a_9929_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X2 a_1993_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X3 a_8937_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X4 w_415_600# a_14135_1380# a_13897_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.72 as=2.975 ps=6.19 w=5 l=0.6
X5 w_415_600# a_3295_1380# a_2985_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X6 a_5961_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X7 w_415_600# a_2303_1380# a_1993_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X8 w_415_600# a_7263_1380# a_6953_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X9 a_4969_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X10 w_415_600# a_11231_1380# a_10921_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X11 a_12905_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X12 w_415_600# a_10239_1380# a_9929_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X13 a_8937_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X14 w_415_600# a_3295_1380# a_2985_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X15 w_415_600# a_2303_1380# a_1993_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X16 w_415_600# a_7263_1380# a_6953_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X17 a_12905_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X18 a_3977_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X19 a_7945_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X20 w_415_600# a_13215_1380# a_12905_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X21 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X22 w_415_600# a_6271_1380# a_5961_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X23 a_3977_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X24 w_415_600# a_5279_1380# a_4969_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X25 a_11913_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X26 a_7945_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X27 a_10921_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X28 w_415_600# a_13215_1380# a_12905_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X29 w_415_600# a_9247_1380# a_8937_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X30 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X31 w_415_600# a_6271_1380# a_5961_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X32 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=4.325 ps=11.73 w=5 l=0.6
X33 w_415_600# a_5279_1380# a_4969_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X34 a_11913_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X35 a_2985_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X36 a_6953_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X37 w_415_600# a_9247_1380# a_8937_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X38 a_10921_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X39 w_415_600# a_12223_1380# a_11913_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X40 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=4.325 ps=11.73 w=5 l=0.6
X41 a_9929_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X42 a_2985_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X43 w_415_600# a_4287_1380# a_3977_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X44 a_6953_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X45 w_415_600# a_8255_1380# a_7945_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X46 w_415_600# a_12223_1380# a_11913_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X47 a_13897_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.975 pd=6.19 as=3.775 ps=11.51 w=5 l=0.6
X48 a_9929_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X49 a_1993_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X50 w_415_600# a_4287_1380# a_3977_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X51 w_415_600# a_14135_1380# a_13897_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.72 as=2.975 ps=6.19 w=5 l=0.6
X52 a_5961_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X53 w_415_600# a_11231_1380# a_10921_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X54 w_415_600# a_8255_1380# a_7945_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X55 a_4969_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
.ends

.subckt sky130_fd_io__top_analog_pad_pudrvr_strong vnb pu_h_n<2> pu_h_n<3> sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_2985_1552#
+ sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_4969_1552# sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_5961_1552#
+ sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_7945_1552# sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/w_415_600#
+ sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_9929_1552# tie_hi_esd sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_11913_1552#
+ sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_1993_1552# sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_13897_1552#
+ sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_3977_1552# a_14575_n152# sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_6953_1552#
+ sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_1001_1552# sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_8937_1552#
+ sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_10921_1552# sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_12905_1552#
Xsky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0 sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/w_415_600#
+ sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_4969_1552# pu_h_n<2> sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_5961_1552#
+ m1_14229_1478# m1_8837_1478# pu_h_n<3> sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_10921_1552#
+ sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_7945_1552# sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_12905_1552#
+ pu_h_n<3> m1_11745_1478# sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_9929_1552#
+ m1_8837_1478# pu_h_n<2> sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_1993_1552#
+ pu_h_n<3> pu_h_n<3> m1_10391_1478# m1_14229_1478# pu_h_n<2> sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_3977_1552#
+ pu_h_n<2> pu_h_n<3> pu_h_n<2> sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_6953_1552#
+ m1_10391_1478# sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_11913_1552#
+ sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_1001_1552# pu_h_n<3> pu_h_n<3>
+ m1_11745_1478# m1_10391_1478# sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_13897_1552#
+ sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_8937_1552# m1_8837_1478# pu_h_n<2>
+ m1_13667_1478# pu_h_n<3> sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad_0/a_2985_1552#
+ m1_11745_1478# pu_h_n<2> pu_h_n<3> sky130_fd_io__PFET_con_diff_wo_abt_270_analog_pad
R0 m2_14075_657# pu_h_n<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X0 tie_hi_esd a_14575_n152# sky130_fd_pr__res_generic_po w=0.5 l=10.2
R1 m1_14229_1478# m2_14532_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 m1_13667_1478# m2_13593_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R3 m2_12849_n185# pu_h_n<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 m1_8837_1478# m2_10673_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 m1_10391_1478# m2_10945_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R6 m2_10673_n208# pu_h_n<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 m2_11422_n209# pu_h_n<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 m1_13667_1478# m2_14075_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 m2_10197_n209# tie_hi_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 m2_10945_n209# tie_hi_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 m1_11745_1478# m2_12608_116# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 m1_10391_1478# m2_11422_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 m1_11745_1478# m2_12849_116# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 m2_12608_n185# pu_h_n<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 m2_13837_658# pu_h_n<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 m2_14769_657# pu_h_n<2> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 m2_11186_n208# pu_h_n<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R18 m2_14286_658# tie_hi_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 m1_8837_1478# m2_10197_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m1_8837_1478# m2_10439_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 m2_14532_657# pu_h_n<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 m1_10391_1478# m2_11186_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R23 m2_13593_657# tie_hi_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 m1_13667_1478# m2_13837_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 m1_14229_1478# m2_14769_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 m1_11745_1478# m2_12365_n184# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 m2_10439_n209# pu_h_n<3> sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 m2_12365_n184# tie_hi_esd sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R29 m1_14229_1478# m2_14286_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__top_analog_pad vccd vddio_q vcchib vssio_q vssd amuxbus_b amuxbus_a
+ pad_core vssa vddio vswitch vdda vssio pad
Xsky130_fd_io__top_analog_pad_pddrvr_strong_0 vssio sky130_fd_io__top_analog_pad_pddrvr_strong_0/pd_h<3>
+ sky130_fd_io__top_analog_pad_pddrvr_strong_0/force_lo_h sky130_fd_io__top_analog_pad_pddrvr_strong_0/pd_h<3>
+ sky130_fd_io__top_analog_pad_pddrvr_strong_0/pd_h<3> sky130_fd_io__top_analog_pad_pddrvr_strong_0/force_lovol_h
+ sky130_fd_io__top_analog_pad_pddrvr_strong_0/vssio_amx vddio pad pad pad pad pad
+ pad pad pad pad pad pad pad vssio pad pad sky130_fd_io__top_analog_pad_pddrvr_strong
Xsky130_fd_io__top_analog_pad_pudrvr_strong_0 vssd sky130_fd_io__top_analog_pad_pudrvr_strong_0/pu_h_n<3>
+ sky130_fd_io__top_analog_pad_pudrvr_strong_0/pu_h_n<3> pad pad pad pad vddio pad
+ sky130_fd_io__top_analog_pad_pudrvr_strong_0/pu_h_n<3> pad pad pad pad vddio pad
+ pad pad pad pad sky130_fd_io__top_analog_pad_pudrvr_strong
R0 pad pad_core sky130_fd_pr__res_generic_m3 w=8.98 l=0.9
.ends

.subckt sky130_fd_io__top_power_lvc_wpad VSSIO_Q VCCHIB VDDA VDDIO_Q P_PAD SRC_BDY_LVC1
+ SRC_BDY_LVC2 BDY2_B2B DRN_LVC2 DRN_LVC1 P_CORE PADISOR PADISOL OGC_LVC AMUXBUS_B
+ VSSIO VDDIO VSSD VSWITCH VSSA AMUXBUS_A VCCD
Xsky130_fd_io__com_busses_esd_0 VCCHIB P_PAD VSSD P_CORE AMUXBUS_A VCCD AMUXBUS_B
+ VDDIO VSSA VSSIO VSWITCH VDDA VDDIO_Q VSSIO_Q sky130_fd_io__com_busses_esd
X0 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X1 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X2 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X3 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X4 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X5 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X6 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X7 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X8 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X9 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X10 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X11 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X12 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X13 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X14 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X15 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X16 SRC_BDY_LVC2 a_2595_15129# a_2872_5340# SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=4.76 ps=15.36 w=7 l=0.18
X17 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X18 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X19 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X20 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X21 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X22 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X23 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X24 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X25 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X26 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X27 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X28 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X29 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X30 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X31 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X32 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X33 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X34 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X35 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X36 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X37 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X38 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X39 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=0 ps=0 w=7 l=8
X40 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X41 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X42 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X43 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X44 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X45 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X46 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.56 w=7 l=0.18
X47 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X48 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X49 a_414_306# DRN_LVC1 sky130_fd_pr__res_generic_po w=0.33 l=1.95k
X50 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X51 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X52 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X53 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X54 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X55 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X56 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X57 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X58 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X59 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X60 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X61 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X62 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X63 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X64 a_2183_16816# a_2595_15129# sky130_fd_pr__res_generic_po w=0.33 l=200
X65 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X66 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X67 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X68 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X69 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X70 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X71 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X72 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X73 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X74 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X75 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X76 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X77 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X78 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X79 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X80 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X81 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X82 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X83 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X84 a_1871_4484# a_13955_3836# sky130_fd_pr__res_generic_po w=0.33 l=300
X85 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X86 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X87 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X88 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X89 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X90 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X91 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X92 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X93 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X94 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X95 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X96 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X97 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X98 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X99 SRC_BDY_LVC1 a_414_306# a_450_404# SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=4.76 ps=15.36 w=7 l=0.18
X100 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X101 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X102 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=0 ps=0 w=7 l=8
X103 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X104 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X105 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X106 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X107 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X108 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X109 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X110 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X111 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X112 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X113 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X114 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X115 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X116 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X117 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X118 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X119 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X120 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X121 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X122 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X123 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X124 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X125 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X126 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X127 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X128 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X129 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X130 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X131 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X132 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X133 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X134 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X135 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X136 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X137 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X138 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X139 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X140 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X141 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=0 ps=0 w=7 l=8
X142 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X143 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X144 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.56 w=7 l=0.18
X145 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X146 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X147 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X148 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X149 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X150 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X151 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X152 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X153 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X154 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X155 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X156 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X157 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X158 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X159 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X160 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X161 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X162 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X163 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X164 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X165 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X166 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X167 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X168 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X169 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X170 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X171 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X172 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X173 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X174 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X175 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X176 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X177 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X178 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X179 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X180 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X181 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X182 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X183 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X184 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X185 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X186 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X187 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X188 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X189 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X190 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X191 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X192 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X193 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X194 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X195 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X196 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X197 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X198 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X199 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X200 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X201 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X202 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X203 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X204 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X205 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X206 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X207 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X208 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X209 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X210 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X211 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X212 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X213 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X214 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X215 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X216 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.56 as=0.98 ps=7.28 w=7 l=0.18
X217 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X218 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X219 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X220 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X221 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X222 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X223 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X224 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X225 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X226 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X227 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X228 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X229 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X230 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X231 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X232 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X233 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X234 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X235 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X236 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X237 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X238 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X239 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X240 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X241 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X242 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X243 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X244 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X245 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X246 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X247 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X248 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X249 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X250 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X251 DRN_LVC2 a_13955_3836# sky130_fd_pr__res_generic_po w=0.33 l=900
X252 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X253 a_1871_4484# a_2183_16816# sky130_fd_pr__res_generic_po w=0.33 l=720
X254 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X255 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X256 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X257 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X258 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X259 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X260 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X261 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.56 as=0.98 ps=7.28 w=7 l=0.18
X262 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X263 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X264 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X265 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X266 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X267 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X268 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X269 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X270 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X271 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X272 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X273 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X274 SRC_BDY_LVC2 a_2595_15129# a_2872_5340# SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=4.76 ps=15.36 w=7 l=0.18
X275 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X276 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X277 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X278 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X279 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X280 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X281 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X282 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X283 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X284 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X285 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=0 ps=0 w=7 l=8
X286 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X287 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X288 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X289 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X290 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X291 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X292 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X293 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X294 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X295 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X296 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X297 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X298 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X299 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X300 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X301 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X302 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X303 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X304 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X305 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X306 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X307 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X308 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X309 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X310 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X311 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X312 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X313 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X314 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X315 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X316 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X317 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X318 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X319 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.56 as=0.98 ps=7.28 w=7 l=0.18
X320 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X321 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X322 SRC_BDY_LVC1 a_414_306# a_450_404# SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=4.76 ps=15.36 w=7 l=0.18
X323 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.56 w=7 l=0.18
X324 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X325 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X326 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X327 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X328 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X329 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X330 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.56 as=0.98 ps=7.28 w=7 l=0.18
X331 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X332 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X333 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X334 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X335 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X336 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X337 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X338 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X339 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X340 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X341 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X342 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X343 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X344 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X345 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X346 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X347 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X348 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X349 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X350 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X351 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X352 SRC_BDY_LVC1 a_414_306# a_450_404# SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=4.76 ps=15.36 w=7 l=0.18
X353 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=0 ps=0 w=7 l=8
X354 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X355 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X356 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X357 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X358 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X359 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X360 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X361 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X362 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X363 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X364 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X365 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X366 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X367 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X368 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X369 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X370 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X371 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X372 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X373 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.56 w=7 l=0.18
X374 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X375 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
R0 P_CORE PADISOL sky130_fd_pr__res_generic_m3 w=12.245 l=10m
X376 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X377 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X378 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X379 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X380 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X381 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X382 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X383 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X384 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X385 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X386 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X387 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X388 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X389 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X390 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X391 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X392 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X393 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X394 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X395 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X396 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X397 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X398 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X399 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X400 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X401 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X402 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X403 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X404 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X405 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X406 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X407 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X408 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X409 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X410 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X411 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X412 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X413 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X414 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X415 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X416 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X417 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X418 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X419 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X420 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X421 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X422 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X423 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X424 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X425 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X426 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X427 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X428 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X429 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X430 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X431 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X432 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X433 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X434 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X435 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X436 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X437 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X438 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X439 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X440 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X441 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X442 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X443 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X444 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=1.325 pd=10.53 as=0 ps=0 w=5 l=4
X445 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X446 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X447 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X448 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X449 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X450 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X451 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X452 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X453 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X454 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X455 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X456 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X457 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X458 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X459 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X460 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X461 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X462 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
R1 P_CORE PADISOR sky130_fd_pr__res_generic_m3 w=12.24 l=10m
X463 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X464 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X465 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
.ends

.subckt sky130_ef_io__vccd_lvc_clamped3_pad VDDA VCCHIB VSSD1 VDDIO AMUXBUS_B VSWITCH
+ VSSIO AMUXBUS_A VCCD VCCD_PAD VCCD1 VSSD VSSA VDDIO_Q VSSIO_Q
Xsky130_fd_io__top_power_lvc_wpad_0 VSSIO_Q VCCHIB VDDA VDDIO_Q VCCD_PAD VSSD1 VSSD1
+ VSSIO VCCD1 VCCD1 VCCD1 sky130_fd_io__top_power_lvc_wpad_0/PADISOR sky130_fd_io__top_power_lvc_wpad_0/PADISOL
+ VSSIO AMUXBUS_B VSSIO VDDIO VSSD VSWITCH VSSA AMUXBUS_A VCCD sky130_fd_io__top_power_lvc_wpad
.ends

.subckt sky130_fd_io__top_ground_lvc_wpad PADISOR PADISOL VSSIO_Q VCCHIB VDDA VDDIO_Q
+ G_PAD SRC_BDY_LVC1 SRC_BDY_LVC2 BDY2_B2B DRN_LVC2 DRN_LVC1 G_CORE OGC_LVC AMUXBUS_B
+ VSSIO VDDIO VSSD VSWITCH VSSA AMUXBUS_A VCCD
Xsky130_fd_io__com_busses_esd_0 VCCHIB G_PAD VSSD G_CORE AMUXBUS_A VCCD AMUXBUS_B
+ VDDIO VSSA VSSIO VSWITCH VDDA VDDIO_Q VSSIO_Q sky130_fd_io__com_busses_esd
X0 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X1 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X2 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X3 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X4 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X5 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X6 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X7 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X8 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X9 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X10 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X11 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X12 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X13 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X14 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X15 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X16 SRC_BDY_LVC2 a_2595_15129# a_2872_5340# SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=4.76 ps=15.36 w=7 l=0.18
X17 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X18 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X19 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X20 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X21 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X22 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X23 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X24 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X25 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X26 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X27 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X28 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X29 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X30 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X31 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X32 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X33 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X34 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X35 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X36 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X37 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X38 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X39 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=0 ps=0 w=7 l=8
X40 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X41 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X42 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X43 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X44 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X45 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X46 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.56 w=7 l=0.18
X47 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X48 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X49 a_414_306# DRN_LVC1 sky130_fd_pr__res_generic_po w=0.33 l=1.95k
X50 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X51 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X52 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X53 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X54 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X55 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X56 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X57 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X58 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X59 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X60 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X61 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X62 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X63 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X64 a_2183_16816# a_2595_15129# sky130_fd_pr__res_generic_po w=0.33 l=200
X65 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X66 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X67 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X68 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X69 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X70 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X71 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X72 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X73 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X74 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X75 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X76 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X77 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X78 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X79 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X80 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X81 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X82 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X83 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X84 a_1871_4484# a_13955_3836# sky130_fd_pr__res_generic_po w=0.33 l=300
X85 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X86 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X87 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X88 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X89 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X90 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X91 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X92 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X93 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X94 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X95 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X96 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X97 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X98 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X99 SRC_BDY_LVC1 a_414_306# a_450_404# SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=4.76 ps=15.36 w=7 l=0.18
X100 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X101 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X102 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=0 ps=0 w=7 l=8
X103 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X104 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X105 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X106 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X107 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X108 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X109 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X110 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X111 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X112 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X113 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X114 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X115 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X116 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X117 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X118 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X119 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X120 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X121 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X122 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X123 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X124 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X125 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X126 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X127 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X128 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X129 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X130 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X131 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X132 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X133 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X134 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X135 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X136 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X137 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X138 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X139 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X140 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X141 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=0 ps=0 w=7 l=8
X142 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X143 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X144 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.56 w=7 l=0.18
X145 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X146 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X147 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X148 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X149 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X150 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X151 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X152 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X153 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X154 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X155 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X156 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X157 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X158 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X159 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X160 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X161 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X162 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X163 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X164 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X165 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X166 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X167 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X168 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X169 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X170 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X171 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X172 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X173 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X174 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X175 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X176 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X177 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X178 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X179 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X180 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X181 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X182 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X183 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X184 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X185 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X186 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X187 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X188 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X189 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X190 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X191 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X192 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X193 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X194 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X195 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X196 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X197 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X198 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X199 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X200 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X201 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X202 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X203 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X204 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X205 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
R0 G_CORE PADISOR sky130_fd_pr__res_generic_m3 w=11.825 l=10m
X206 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X207 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X208 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X209 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X210 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X211 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X212 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X213 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X214 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X215 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X216 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.56 as=0.98 ps=7.28 w=7 l=0.18
X217 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X218 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X219 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X220 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X221 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X222 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X223 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X224 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X225 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X226 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
R1 G_CORE PADISOL sky130_fd_pr__res_generic_m3 w=11.825 l=10m
X227 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X228 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X229 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X230 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X231 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X232 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X233 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X234 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X235 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X236 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X237 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X238 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X239 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X240 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X241 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X242 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X243 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X244 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X245 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X246 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X247 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X248 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X249 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X250 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X251 DRN_LVC2 a_13955_3836# sky130_fd_pr__res_generic_po w=0.33 l=900
X252 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X253 a_1871_4484# a_2183_16816# sky130_fd_pr__res_generic_po w=0.33 l=720
X254 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X255 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X256 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X257 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X258 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X259 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X260 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X261 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.56 as=0.98 ps=7.28 w=7 l=0.18
X262 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X263 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X264 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X265 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X266 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X267 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X268 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X269 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X270 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X271 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X272 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X273 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X274 SRC_BDY_LVC2 a_2595_15129# a_2872_5340# SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=4.76 ps=15.36 w=7 l=0.18
X275 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X276 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X277 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X278 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X279 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X280 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X281 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X282 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X283 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X284 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X285 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=0 ps=0 w=7 l=8
X286 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X287 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X288 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X289 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X290 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X291 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X292 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X293 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X294 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X295 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X296 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X297 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X298 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X299 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X300 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X301 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X302 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X303 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X304 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X305 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X306 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X307 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X308 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X309 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X310 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X311 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X312 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X313 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X314 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X315 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X316 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X317 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X318 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X319 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.56 as=0.98 ps=7.28 w=7 l=0.18
X320 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X321 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X322 SRC_BDY_LVC1 a_414_306# a_450_404# SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=4.76 ps=15.36 w=7 l=0.18
X323 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.56 w=7 l=0.18
X324 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X325 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X326 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X327 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X328 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X329 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X330 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.56 as=0.98 ps=7.28 w=7 l=0.18
X331 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X332 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X333 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X334 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X335 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X336 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X337 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X338 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X339 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X340 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X341 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X342 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X343 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X344 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X345 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X346 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X347 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X348 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X349 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X350 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X351 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X352 SRC_BDY_LVC1 a_414_306# a_450_404# SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=4.76 ps=15.36 w=7 l=0.18
X353 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.3975 pd=7.685 as=0 ps=0 w=7 l=8
X354 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X355 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X356 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X357 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X358 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X359 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X360 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X361 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X362 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X363 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X364 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X365 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X366 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X367 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X368 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X369 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X370 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X371 SRC_BDY_LVC1 BDY2_B2B sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X372 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X373 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.56 w=7 l=0.18
X374 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X375 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X376 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X377 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X378 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X379 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X380 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X381 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X382 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X383 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X384 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X385 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X386 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X387 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X388 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X389 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X390 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X391 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X392 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X393 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X394 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X395 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X396 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X397 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X398 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X399 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X400 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X401 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X402 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X403 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X404 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X405 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X406 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X407 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=5.625 pd=12.25 as=2.925 ps=6.17 w=5 l=0.18
X408 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X409 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X410 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X411 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X412 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X413 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X414 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X415 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X416 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X417 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X418 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X419 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X420 SRC_BDY_LVC1 a_414_306# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X421 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X422 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X423 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X424 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X425 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X426 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X427 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X428 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X429 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X430 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X431 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X432 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X433 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X434 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X435 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X436 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X437 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X438 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X439 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X440 BDY2_B2B SRC_BDY_LVC1 sky130_fd_pr__diode_pd2nw_05v5 perim=3.3e+07 area=2.25e+13
X441 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X442 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X443 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X444 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=1.325 pd=10.53 as=0 ps=0 w=5 l=4
X445 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X446 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X447 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X448 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X449 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X450 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
X451 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X452 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X453 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X454 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X455 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=6.17 as=5.625 ps=12.25 w=5 l=0.18
X456 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X457 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X458 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.535 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X459 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.525 ps=6.01 w=5 l=0.18
X460 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X461 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=7.875 pd=16.25 as=4.095 ps=8.17 w=7 l=0.18
X462 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X463 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.525 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X464 SRC_BDY_LVC1 a_450_404# DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.535 ps=8.01 w=7 l=0.18
X465 DRN_LVC1 a_450_404# SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 ad=4.095 pd=8.17 as=7.875 ps=16.25 w=7 l=0.18
.ends

.subckt sky130_ef_io__vssd_lvc_clamped3_pad VDDA VSSIO_Q VSSD1 VCCD VSSD VSSA AMUXBUS_B
+ AMUXBUS_A VSSD_PAD VSWITCH VDDIO VCCHIB VDDIO_Q VSSIO VCCD1
Xsky130_fd_io__top_ground_lvc_wpad_1 sky130_fd_io__top_ground_lvc_wpad_1/PADISOR sky130_fd_io__top_ground_lvc_wpad_1/PADISOL
+ VSSIO_Q VCCHIB VDDA VDDIO_Q VSSD_PAD VSSD1 VSSD1 VSSIO VCCD1 VCCD1 VSSD1 VSSIO AMUXBUS_B
+ VSSIO VDDIO VSSD VSWITCH VSSA AMUXBUS_A VCCD sky130_fd_io__top_ground_lvc_wpad
.ends

* Black-box entry subcircuit for sky130_fd_io__top_sio_macro abstract view
.subckt sky130_fd_io__top_sio_macro vssa vddio vccd vcchib vdda vddio_q vssd vssio
+ vswitch vssio_q pad<1> pad<0> amuxbus_b amuxbus_a vreg_en_refgen hld_h_n_refgen
+ voh_sel<0> voh_sel<1> voh_sel<2> vohref enable_vdda_h vtrip_sel_refgen dft_refgen
+ dm1<1> dm1<2> dm1<0> dm0<0> dm0<1> dm0<2> voutref_dft ibuf_sel_refgen vref_sel<0>
+ pad_a_esd_1_h<0> ibuf_sel<1> vinref_dft pad_a_esd_1_h<1> pad_a_esd_0_h<1> vref_sel<1>
+ pad_a_esd_0_h<0> pad_a_noesd_h<0> pad_a_noesd_h<1> inp_dis<1> inp_dis<0> tie_lo_esd<0>
+ tie_lo_esd<1> out<1> out<0> vtrip_sel<0> vtrip_sel<1> enable_h vreg_en<0> vreg_en<1>
+ slow<1> slow<0> oe_n<0> oe_n<1> in_h<1> in_h<0> in<0> in<1> hld_ovr<1> hld_ovr<0>
+ hld_h_n<1> hld_h_n<0> ibuf_sel<0>
.ends

.subckt sky130_fd_io__top_vrefcapv2 cpos cneg vssio vddio_q vddio vssio_q vccd vssa
+ vcchib vswitch vdda vssd amuxbus_b amuxbus_a
X0 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X1 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X2 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X3 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X4 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X5 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X6 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X7 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X8 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X9 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X10 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X11 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X12 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X13 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X14 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X15 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X16 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X17 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X18 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X19 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X20 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X21 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X22 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X23 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X24 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X25 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X26 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X27 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X28 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X29 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X30 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X31 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X32 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X33 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X34 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X35 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X36 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X37 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X38 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X39 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X40 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X41 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X42 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X43 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X44 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X45 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X46 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X47 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X48 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X49 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X50 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X51 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X52 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X53 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X54 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X55 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X56 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X57 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X58 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X59 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X60 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X61 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X62 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X63 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X64 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X65 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X66 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X67 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X68 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X69 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X70 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X71 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X72 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X73 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X74 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X75 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X76 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X77 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X78 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X79 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X80 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X81 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X82 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X83 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X84 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X85 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X86 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X87 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X88 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X89 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X90 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X91 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X92 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X93 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X94 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X95 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X96 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X97 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X98 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X99 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X100 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X101 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X102 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X103 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X104 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X105 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X106 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X107 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X108 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X109 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X110 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X111 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X112 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X113 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X114 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X115 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X116 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X117 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X118 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X119 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X120 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X121 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X122 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X123 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X124 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X125 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X126 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X127 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X128 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X129 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X130 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X131 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X132 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X133 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X134 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X135 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X136 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X137 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X138 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X139 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X140 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X141 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X142 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X143 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X144 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X145 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X146 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X147 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X148 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X149 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X150 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X151 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X152 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X153 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X154 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X155 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X156 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X157 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X158 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X159 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X160 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X161 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=0.9
X162 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X163 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X164 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X165 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X166 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X167 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X168 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X169 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X170 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X171 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X172 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X173 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X174 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X175 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X176 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X177 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X178 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
X179 cneg cpos cneg cneg sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=0.9
.ends

.subckt sky130_ef_io__vdda_hvc_clamped_pad VDDIO_Q VSSIO_Q VSSIO VDDA_PAD AMUXBUS_B
+ AMUXBUS_A VDDA VSSD VCCHIB VSSA VDDIO VSWITCH VCCD
Xsky130_fd_io__top_power_hvc_wpadv2_1 VSSA VDDIO AMUXBUS_B VDDA VSSIO_Q VDDA_PAD sky130_fd_io__top_power_hvc_wpadv2_1/PADISOL
+ VDDIO_Q VDDA sky130_fd_io__top_power_hvc_wpadv2_1/PADISOR VDDA VCCHIB VCCD VSWITCH
+ VDDIO VSSA VSSD AMUXBUS_A VSSIO sky130_fd_io__top_power_hvc_wpadv2
.ends

.subckt sky130_fd_io__com_res_weak_v2 a_n281_1306# a_534_6146#
X0 a_n281_1656# a_n281_1306# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R0 a_n13_3671# m1_3_3617# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X1 a_n283_3382# a_n283_2797# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R1 m1_n268_3094# a_n283_2797# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R2 m1_n268_1364# a_n281_1306# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R3 m1_3_3580# a_n13_2329# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X2 a_n283_2797# a_n283_2447# sky130_fd_pr__res_generic_po w=0.8 l=1.5
X3 a_n13_3671# a_n13_2329# sky130_fd_pr__res_generic_po w=0.8 l=6
R4 a_n283_2447# m1_n268_1924# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R5 a_n283_2797# m1_n268_2513# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
X4 a_n13_2329# a_n283_3382# sky130_fd_pr__res_generic_po w=0.8 l=6
R6 a_n13_2329# m1_2_2233# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R7 m1_n268_1924# a_n281_1656# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
X5 a_n13_6243# a_534_6146# sky130_fd_pr__res_generic_po w=0.8 l=50
X6 a_n13_6243# a_n13_3671# sky130_fd_pr__res_generic_po w=0.8 l=12
R8 m1_n268_2513# a_n283_2447# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R9 m1_2_2233# a_n283_3382# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X7 a_n283_2447# a_n281_1656# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R10 a_n283_3382# m1_n268_3094# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R11 a_n281_1656# m1_n268_1364# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
.ends

.subckt sky130_fd_io__xres4v2_in_buf VGND IN_H VDDIO VNORMAL VNORMAL_B PAD ENABLE_HV
+ IN_H_N VCCHIB ENABLE_VDDIO_LV a_n445_2580# m2_288_2575# w_4058_2188# a_n32352_n9635#
Xsky130_fd_io__inv_1_0 VGND VCCHIB VCCHIB VGND sky130_fd_io__inv_1_0/Y ENABLE_VDDIO_LV
+ sky130_fd_io__inv_1
X0 a_n29280_n8739# VNORMAL_B a_n31524_n8739# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.56 w=5 l=0.5
X1 a_n11573_n8777# a_111_449# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X2 VGND a_n176_869# a_2300_3398# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X3 a_1560_2580# ENABLE_HV VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.795 ps=6.53 w=3 l=0.5
X4 VGND IN_H_N IN_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X5 VGND PAD a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X6 a_n232_901# a_n176_869# a_469_2037# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.56 as=0.7 ps=5.28 w=5 l=0.8
X7 a_2165_2545# a_n176_869# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.795 ps=6.53 w=3 l=0.5
X8 VGND a_2165_2545# a_2356_3115# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X9 VDDIO a_2356_3115# a_2300_3398# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.5
X10 IN_H_N a_2300_3398# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.795 ps=6.53 w=3 l=0.5
X11 a_5826_2675# ENABLE_HV VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X12 a_n176_869# PAD w_5030_2188# w_5030_2188# sky130_fd_pr__pfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=0.8
X13 a_n16_901# a_n176_869# a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.56 as=1.4 ps=10.56 w=5 l=0.8
X14 a_1560_2580# ENABLE_HV VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.56 as=1.325 ps=10.53 w=5 l=0.5
X15 a_n232_901# PAD VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X16 IN_H IN_H_N VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.42 ps=3.28 w=3 l=0.5
X17 VDDIO a_5826_2675# a_111_449# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X18 IN_H_N a_2300_3398# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.795 ps=6.53 w=3 l=0.5
X19 VGND a_5826_2675# a_111_449# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.1855 ps=1.93 w=0.7 l=0.6
X20 a_2356_3115# a_2165_2545# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X21 VDDIO a_111_449# a_n29280_n8739# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X22 VDDIO VNORMAL_B a_5826_2675# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X23 a_n176_869# PAD a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.56 w=5 l=0.8
X24 a_n9813_4210# VNORMAL_B a_n11573_n8777# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X25 VGND VNORMAL_B a_5852_3096# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X26 a_2300_3398# a_n176_869# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X27 w_4058_2188# a_111_449# a_n445_2580# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=0.9
X28 VGND VGND VGND VGND sky130_fd_pr__nfet_05v0_nvt ad=2.65 pd=20.53 as=0 ps=0 w=10 l=0.9
X29 a_2165_2545# a_n176_869# w_4058_2188# w_4058_2188# sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.56 as=1.4 ps=10.56 w=5 l=0.5
X30 IN_H IN_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.5
X31 IN_H IN_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X32 a_469_2037# a_n176_869# a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X33 VDDIO IN_H_N IN_H VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X34 a_n757_2580# a_111_449# w_5030_2188# VGND sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=2.8 ps=20.56 w=10 l=0.9
X35 a_n16_901# VNORMAL_B VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.56 as=0.7 ps=5.28 w=5 l=0.5
X36 a_n232_901# PAD a_n176_869# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X37 a_n29280_n8739# a_n31524_n8739# VGND sky130_fd_pr__res_generic_nd__hv w=0.29 l=1.07719k
X38 VCCHIB sky130_fd_io__inv_1_0/Y a_n757_2580# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.56 w=5 l=0.5
X39 w_5030_2188# w_5030_2188# w_5030_2188# w_5030_2188# sky130_fd_pr__pfet_g5v0d10v5 ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.8
X40 a_n232_901# a_n176_869# a_469_2037# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X41 a_5826_2675# ENABLE_HV VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X42 VDDIO a_5826_2675# a_111_449# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X43 a_n176_869# PAD a_n31524_n8739# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.56 as=1.4 ps=10.56 w=5 l=0.5
X44 a_2165_2545# a_n176_869# a_n9813_4210# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.56 as=0.7 ps=5.28 w=5 l=0.5
X45 a_469_2037# PAD a_157_2580# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=0.9
X46 a_5852_3096# ENABLE_HV a_5826_2675# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X47 a_n9813_4210# a_n11573_n8777# sky130_fd_pr__res_generic_po w=0.4 l=713.69501
X48 IN_H IN_H_N VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X49 VDDIO VNORMAL_B a_5826_2675# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X50 a_2356_3115# a_2300_3398# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1176 pd=1.4 as=0.0588 ps=0.7 w=0.42 l=0.5
X51 a_n445_2580# sky130_fd_io__inv_1_0/Y VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.56 as=0.7 ps=5.28 w=5 l=0.5
X52 VDDIO VNORMAL a_157_2580# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.56 w=5 l=0.5
X53 a_469_2037# a_n176_869# a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
.ends

.subckt sky130_fd_io__xres_inv_hysv2 VCC_IO VSSD OUT_H a_122_112# a_322_144# a_322_604#
X0 a_322_144# OUT_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1176 pd=1.4 as=0.1176 ps=1.4 w=0.42 l=1
X1 a_578_144# a_122_112# a_322_604# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.42 ps=3.28 w=3 l=1
X2 a_322_144# a_122_112# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=1
X3 a_578_144# a_122_112# a_322_144# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=1
X4 OUT_H a_578_144# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X5 VCC_IO OUT_H a_322_604# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.1176 pd=1.4 as=0.1176 ps=1.4 w=0.42 l=1
X6 OUT_H a_578_144# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=0.5
X7 a_322_604# a_122_112# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.84 ps=6.56 w=3 l=1
.ends

.subckt sky130_fd_io__gpio_buf_localesdv2 VTRIP_SEL_H OUT_H OUT_VT sky130_fd_io__res250only_small_0/PAD
+ VGND VCC_IO
Xsky130_fd_io__signal_5_sym_hv_local_5term_0 VGND VCC_IO OUT_VT VGND VCC_IO VCC_IO
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_1 VGND VCC_IO VGND VGND OUT_VT VCC_IO sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_2 VGND VCC_IO OUT_H VGND VCC_IO VCC_IO
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_3 VGND VCC_IO VGND VGND OUT_H VCC_IO sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__res250only_small_0 sky130_fd_io__res250only_small_0/PAD OUT_H sky130_fd_io__res250only_small
X0 OUT_VT VTRIP_SEL_H OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=1
.ends

.subckt sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2 VCC_IO a_10282_1285# a_5322_1285#
+ a_8980_1457# a_7988_1457# a_2036_1457# a_13940_1457# a_12948_1457# a_12266_1285#
+ a_7306_1285# a_5012_1457# a_3900_1285# a_2908_1285# a_5884_1285# a_14178_1285# a_10844_1285#
+ a_1354_1285# a_7868_1285# a_12828_1285# a_8860_1285# a_13820_1285# a_4330_1285#
+ a_3338_1285# a_6996_1457# a_11956_1457# a_1044_1457# a_11274_1285# a_6314_1285#
+ w_469_785# a_9972_1457# a_4020_1457# a_3028_1457# a_8298_1285# a_13258_1285# a_9290_1285#
+ a_1916_1285# a_6004_1457# a_4892_1285# a_6876_1285# a_924_1285# a_11836_1285# a_2346_1285#
+ a_9852_1285# a_10964_1457#
X0 a_10964_1457# a_10844_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X1 a_9972_1457# a_9852_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X2 w_469_785# a_2346_1285# a_2036_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X3 a_2036_1457# a_1916_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X4 a_6996_1457# a_6876_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X5 w_469_785# a_12266_1285# a_11956_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X6 w_469_785# a_6314_1285# a_6004_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X7 a_11956_1457# a_11836_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X8 w_469_785# a_9290_1285# a_8980_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X9 a_5012_1457# a_4892_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X10 w_469_785# a_4330_1285# a_4020_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X11 a_8980_1457# a_8860_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X12 w_469_785# a_10282_1285# a_9972_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X13 w_469_785# a_3338_1285# a_3028_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X14 w_469_785# a_8298_1285# a_7988_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X15 a_1044_1457# a_924_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.425 ps=11.37 w=5 l=0.6
X16 a_4020_1457# a_3900_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X17 a_13940_1457# a_13820_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=2.975 pd=6.19 as=3.775 ps=11.51 w=5 l=0.6
X18 a_3028_1457# a_2908_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X19 a_7988_1457# a_7868_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X20 w_469_785# a_13258_1285# a_12948_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X21 w_469_785# a_7306_1285# a_6996_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X22 a_12948_1457# a_12828_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X23 w_469_785# a_14178_1285# a_13940_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.425 pd=11.37 as=2.975 ps=6.19 w=5 l=0.6
X24 w_469_785# a_1354_1285# a_1044_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X25 a_6004_1457# a_5884_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X26 w_469_785# a_11274_1285# a_10964_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X27 w_469_785# a_5322_1285# a_5012_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X28 a_9972_1457# a_9852_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X29 a_10964_1457# a_10844_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X30 w_469_785# a_2346_1285# a_2036_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X31 a_6996_1457# a_6876_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X32 w_469_785# a_6314_1285# a_6004_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X33 a_2036_1457# a_1916_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X34 w_469_785# a_12266_1285# a_11956_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X35 a_11956_1457# a_11836_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X36 a_5012_1457# a_4892_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X37 w_469_785# a_9290_1285# a_8980_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X38 a_8980_1457# a_8860_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X39 w_469_785# a_10282_1285# a_9972_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X40 w_469_785# a_4330_1285# a_4020_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X41 a_1044_1457# a_924_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.425 ps=11.37 w=5 l=0.6
X42 a_4020_1457# a_3900_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X43 w_469_785# a_3338_1285# a_3028_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X44 w_469_785# a_8298_1285# a_7988_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X45 a_3028_1457# a_2908_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X46 a_7988_1457# a_7868_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X47 w_469_785# a_7306_1285# a_6996_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X48 a_13940_1457# a_13820_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=2.975 pd=6.19 as=3.775 ps=11.51 w=5 l=0.6
X49 w_469_785# a_13258_1285# a_12948_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X50 a_12948_1457# a_12828_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X51 w_469_785# a_1354_1285# a_1044_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X52 w_469_785# a_14178_1285# a_13940_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.425 pd=11.37 as=2.975 ps=6.19 w=5 l=0.6
X53 a_6004_1457# a_5884_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X54 w_469_785# a_5322_1285# a_5012_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X55 w_469_785# a_11274_1285# a_10964_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpio_pddrvr_strong_xres4v2 PD_H[2] PD_H[3] TIE_LO_ESD VGND_IO
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_11956_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_6996_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_1044_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_9972_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_3028_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_4020_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_6004_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_10964_1457#
+ w_335_3259# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_12948_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_7988_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_13940_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_8980_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_2036_1457# m1_785_3898# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_5012_1457#
+ VCC_IO
Xsky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0 VCC_IO PD_H[3] m1_9769_3903# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_8980_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_7988_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_2036_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_13940_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_12948_1457#
+ m1_2697_3903# m1_7657_3903# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_5012_1457#
+ m1_11193_3903# m1_11193_3903# m1_8232_3903# m1_785_3898# PD_H[3] m1_12747_3903#
+ PD_H[2] m1_2135_3903# PD_H[2] m1_785_3898# m1_9769_3903# m1_11193_3903# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_6996_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_11956_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_1044_1457#
+ PD_H[3] m1_8232_3903# w_335_3259# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_9972_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_4020_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_3028_1457#
+ PD_H[2] m1_785_3898# PD_H[3] m1_12747_3903# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_6004_1457#
+ m1_9769_3903# m1_8232_3903# m1_12747_3903# PD_H[3] m1_12747_3903# PD_H[3] sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_10964_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2
R0 m1_2697_3903# m2_2790_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R1 m2_12763_1099# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 m2_6804_1099# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R3 m1_2135_3903# m2_1848_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 m2_13622_1100# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 m1_12747_3903# m2_12763_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R6 m2_1260_1100# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 m1_7657_3903# m2_6804_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 m2_897_1099# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 m1_12747_3903# m2_13622_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 m1_2135_3903# m2_1260_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 m1_785_3898# m2_897_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 m2_12189_1099# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 m2_9986_1099# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 m2_413_1100# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 m2_3095_1099# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 m2_9366_1099# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 m1_11193_3903# m2_12189_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R18 m1_2697_3903# m2_3095_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 m1_9769_3903# m2_9986_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m1_785_3898# m2_413_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 m1_8232_3903# m2_9366_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 m2_11758_1100# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R23 m1_11193_3903# m2_11758_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 m2_8935_1100# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 m2_10846_1099# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 m2_11329_1099# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 m2_656_1099# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 m2_1565_1099# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R29 m2_3378_1099# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R30 m1_8232_3903# m2_8935_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R31 m1_9769_3903# m2_10846_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R32 m1_11193_3903# m2_11329_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R33 m2_8506_1099# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R34 m2_10415_1100# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R35 m1_785_3898# m2_656_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R36 m2_7664_1099# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R37 m1_2135_3903# m2_1565_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R38 m1_2697_3903# m2_3378_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R39 m1_8232_3903# m2_8506_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R40 m1_9769_3903# m2_10415_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R41 m1_7657_3903# m2_7664_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R42 m2_7233_1100# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R43 m2_13193_1099# PD_H[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R44 m2_2790_1100# PD_H[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R45 m1_7657_3903# m2_7233_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R46 m1_12747_3903# m2_13193_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X0 TIE_LO_ESD VGND_IO sky130_fd_pr__res_generic_po w=0.5 l=10.2
R47 m2_1848_1099# TIE_LO_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__tk_tie_r_out_esd A B
X0 A B sky130_fd_pr__res_generic_po w=0.5 l=10.2
.ends

.subckt sky130_fd_io__xres2v2_rcfilter_lpfv2 IN VCC_IO a_9105_2295# a_1381_4189# a_7373_4189#
+ a_3949_4189# a_2237_4189# a_525_4189# a_472_471# a_7393_2295# a_472_1087# a_8249_2295#
+ a_5661_4189# a_472_779# a_336_26# a_472_317# a_472_1549# a_6517_4189# a_6537_2295#
+ a_9941_4189# a_472_163# a_3093_4189# a_472_1395# a_4805_4189# a_9961_2295# a_9085_4189#
+ a_472_1857#
R0 a_472_1857# m1_3338_1932# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R1 m1_3363_1420# a_3382_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R2 a_472_1087# m1_467_1076# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R3 a_11618_3687# m1_14484_3916# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X0 a_472_7036# a_472_7036# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R4 m1_467_1355# a_472_317# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R5 a_7373_4189# m1_11612_5169# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X1 a_472_1087# a_3382_1087# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R6 m1_14480_3712# a_11618_3687# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R7 m1_467_740# a_472_317# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X2 VCC_IO a_2237_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R8 m1_3363_188# a_3382_163# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R9 a_6517_4189# m1_14484_5691# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R10 a_11618_2147# m1_14484_2376# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X3 a_3382_1703# a_11618_2147# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R11 a_11618_3071# m1_14484_3300# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R12 m1_14480_4922# a_7373_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R13 m1_14480_2172# a_11618_2147# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R14 IN m1_14484_4202# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R15 m1_11613_5471# a_7373_4189# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R16 m1_14328_5846# a_5661_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X4 a_472_6420# a_472_6420# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X5 a_472_6112# a_12884_6112# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X6 a_472_779# a_3382_779# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R17 a_472_6420# m1_3338_6444# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R18 m1_14480_5846# a_5661_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R19 m1_3363_1728# a_3382_1703# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R20 m1_14480_3096# a_11618_3071# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R21 a_7373_4189# m1_14484_5126# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R22 a_472_317# m1_3338_341# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X7 a_472_7344# a_472_7344# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X8 a_472_7036# a_12884_7036# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R23 a_472_7344# m1_3338_7368# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R24 a_472_1395# m1_467_1384# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X9 a_472_317# a_7393_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R25 a_472_779# m1_467_769# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X10 a_472_1395# a_3382_1395# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R26 m1_3334_1112# a_472_1087# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R27 a_472_1857# m1_5939_1932# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X11 a_3382_1087# a_11618_2763# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R28 m1_3363_496# a_3382_471# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X12 a_11618_2147# a_12884_1857# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R29 a_11618_2455# m1_14484_2684# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R30 a_472_1395# m1_10927_1419# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X13 VCC_IO a_7373_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R31 a_472_6728# m1_3338_6752# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X14 a_472_6420# a_12884_6420# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R32 a_472_317# m1_5624_734# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X15 a_472_7652# a_472_7652# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R33 a_7373_4189# m1_14484_5434# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X16 a_472_7344# a_12884_7344# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R34 a_472_7652# m1_3338_7676# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X17 a_472_163# a_3382_163# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R35 a_472_317# m1_6480_426# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X18 a_3382_1395# a_11618_2455# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X19 a_472_317# a_8249_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X20 a_11618_2455# a_12884_1549# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R36 m1_3363_1112# a_3382_1087# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R37 a_11618_2763# m1_14484_2992# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R38 m1_14299_5846# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X21 a_11618_3379# a_12884_625# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R39 m1_467_432# a_472_317# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R40 a_472_317# m1_4825_1042# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R41 a_472_317# m1_6537_426# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X22 a_7373_4189# a_12884_6728# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R42 a_472_317# m1_4768_1042# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R43 a_6517_4189# m1_14484_5742# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X23 a_472_7652# a_12884_7652# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X24 VCC_IO a_7373_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X25 a_9085_4189# a_12884_7344# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X26 a_472_471# a_3382_471# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X27 a_11618_2763# a_12884_1241# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R44 a_472_7036# m1_3338_7060# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R45 a_472_471# m1_467_461# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X28 a_11618_3687# a_12884_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R46 a_472_7344# m1_3338_7419# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X29 a_3382_779# a_11618_3071# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R47 m1_2201_1652# a_472_1549# sky130_fd_pr__res_generic_m1 w=0.29 l=10m
X30 a_6517_4189# a_12884_6420# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X31 a_472_317# a_472_779# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R48 a_472_317# m1_3338_700# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X32 a_7373_4189# a_12884_7036# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R49 m1_10929_804# a_472_779# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X33 a_472_317# a_472_471# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X34 a_472_317# a_472_1857# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X35 a_472_1549# a_472_1549# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R50 a_472_6728# m1_3338_6803# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R51 a_7373_4189# m1_11741_5169# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R52 a_472_7652# m1_3338_7727# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R53 a_472_317# m1_2201_1681# sky130_fd_pr__res_generic_m1 w=0.29 l=10m
X36 VCC_IO a_5661_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R54 m1_10929_188# a_472_163# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X37 VCC_IO a_3949_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X38 a_5661_4189# a_12884_6112# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X39 a_11618_3071# a_12884_933# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R55 a_472_1549# m1_466_1664# sky130_fd_pr__res_generic_m1 w=0.29 l=0.31
R56 a_472_6112# m1_3338_6187# sky130_fd_pr__res_generic_m1 w=0.29 l=0.31
X40 a_472_7652# a_3382_7806# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X41 a_3382_163# a_11618_3687# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X42 a_472_317# a_472_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R57 m1_3334_6907# a_472_6728# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X43 a_472_317# a_6537_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X44 a_472_1857# a_472_1857# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X45 a_472_1549# a_12884_1549# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X46 a_9941_4189# a_12884_7652# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X47 a_11618_2455# a_11618_2455# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X48 a_472_6112# a_3382_6266# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R58 m1_10929_496# a_472_471# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R59 a_472_7036# m1_3338_7111# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X49 VCC_IO a_6517_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X50 a_3382_7806# IN a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X51 a_3382_471# a_11618_3379# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R60 a_472_6420# m1_3338_6495# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R61 a_472_317# m1_3338_392# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X52 a_472_317# a_472_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X53 a_472_1857# a_12884_1857# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R62 m1_3363_6907# a_3382_6882# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X54 a_11618_2763# a_11618_2763# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R63 a_11618_2147# m1_14484_2325# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X55 a_472_317# a_9105_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X56 a_472_6420# a_3382_6574# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X57 a_3382_6266# a_6517_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X58 a_472_317# a_472_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R64 m1_10958_804# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R65 a_11618_3071# m1_14484_3249# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X59 a_472_317# a_472_1549# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=1.855 pd=14.53 as=0 ps=0 w=7 l=4
R66 m1_3334_7215# a_472_7036# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R67 a_472_317# m1_3338_1265# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X60 a_472_7344# a_3382_7498# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X61 a_472_317# a_472_1395# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R68 a_472_1395# m1_10927_1470# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R69 m1_3334_6599# a_472_6420# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R70 a_472_317# m1_3113_1350# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R71 a_9941_4189# m1_14484_4459# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X62 a_472_317# a_472_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R72 a_472_317# m1_3056_1350# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X63 VCC_IO a_3093_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R73 m1_10958_188# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X64 VCC_IO a_525_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.855 pd=14.53 as=0 ps=0 w=7 l=4
R74 a_11618_2455# m1_14484_2633# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X65 IN IN a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X66 a_472_6728# a_3382_6882# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R75 a_11618_3379# m1_14484_3557# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X67 a_3382_6574# a_7373_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X68 a_472_317# a_12884_1241# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R76 a_472_1549# m1_3338_1573# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X69 a_11618_2147# a_11618_2147# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R77 m1_3334_7523# a_472_7344# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R78 a_5661_4189# m1_11613_5808# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X70 a_3382_7498# a_9941_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R79 m1_3363_7215# a_3382_7190# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R80 m1_14509_2480# a_12884_1549# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X71 a_11618_3071# a_11618_3071# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R81 m1_3363_6599# a_3382_6574# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R82 m1_10929_1728# a_472_1549# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R83 a_9085_4189# m1_14484_4767# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X72 a_472_317# a_12884_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R84 m1_14509_4306# a_12884_7652# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R85 m1_3334_804# a_472_779# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R86 a_472_317# m1_3338_1008# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X73 a_472_317# a_472_163# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R87 m1_10958_496# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R88 m1_11613_4547# a_9941_4189# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R89 m1_14509_5230# a_12884_6728# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X74 a_9941_4189# a_9941_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R90 m1_1345_1960# a_472_1857# sky130_fd_pr__res_generic_m1 w=0.29 l=10m
R91 a_11618_2763# m1_14484_2941# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X75 a_3382_6882# a_7373_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X76 a_7373_4189# a_7373_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R92 a_472_1857# m1_3338_1881# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R93 a_11618_3687# m1_14484_3865# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R94 m1_3334_7831# a_472_7652# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R95 m1_14509_3404# a_12884_625# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X77 VCC_IO a_4805_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R96 m1_3363_7523# a_3382_7498# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R97 m1_3334_188# a_472_163# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R98 m1_14509_2788# a_12884_1241# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X78 a_11618_3379# a_11618_3379# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R99 a_472_1549# m1_595_1664# sky130_fd_pr__res_generic_m1 w=0.29 l=0.31
X79 a_472_7036# a_3382_7190# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R100 m1_14509_4614# a_12884_7344# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X80 a_472_317# a_12884_625# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R101 m1_3334_6291# a_472_6112# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R102 a_472_317# m1_3338_1316# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R103 m1_10958_1728# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R104 a_9085_4189# m1_11613_4576# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R105 a_472_317# m1_1345_1989# sky130_fd_pr__res_generic_m1 w=0.29 l=10m
X81 a_9085_4189# a_9085_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R106 m1_10929_1112# a_472_1087# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R107 IN m1_14484_4151# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R108 m1_11613_4855# a_9085_4189# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R109 m1_14509_5538# a_12884_6420# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X82 a_6517_4189# a_6517_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R110 m1_14480_2480# a_11618_2455# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R111 a_9941_4189# m1_14484_4510# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R112 a_7373_4189# m1_14484_5075# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R113 m1_11613_5779# a_6517_4189# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X83 a_472_6728# a_472_6728# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X84 a_472_317# a_9961_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R114 m1_14509_3712# a_12884_317# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R115 a_472_317# m1_3338_649# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R116 m1_3363_7831# a_3382_7806# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R117 m1_14480_4306# a_9941_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R118 a_472_1857# m1_5939_1881# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X85 a_11618_3687# a_11618_3687# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R119 m1_3334_496# a_472_471# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X86 VCC_IO a_9085_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R120 m1_3334_1420# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R121 m1_14480_5230# a_7373_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R122 a_11618_3379# m1_14484_3608# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R123 a_6517_4189# m1_11613_5500# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X87 a_3382_7190# a_9085_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X88 VCC_IO a_1381_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
X89 a_472_317# a_12884_933# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R124 a_472_1549# m1_3338_1624# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R125 m1_14509_2172# a_12884_1857# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R126 m1_14509_4922# a_12884_7036# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R127 m1_467_1047# a_472_317# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R128 a_7373_4189# m1_11613_4884# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X90 VCC_IO a_9941_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R129 m1_3363_6291# a_3382_6266# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R130 m1_14480_3404# a_11618_3379# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R131 m1_14509_5846# a_12884_6112# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R132 a_472_317# m1_5681_734# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R133 m1_14509_3096# a_12884_933# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R134 m1_10958_1112# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R135 m1_14480_2788# a_11618_2763# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R136 a_9085_4189# m1_14484_4818# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R137 a_7373_4189# m1_14484_5383# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X91 a_472_6728# a_12884_6728# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X92 a_472_1549# a_3382_1703# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X93 a_472_317# a_472_1087# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=4
R138 m1_14480_4614# a_9085_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R139 m1_3363_804# a_3382_779# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R140 a_472_317# m1_3338_957# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X94 a_472_6112# a_472_6112# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X95 a_7373_4189# a_7373_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R141 m1_3334_1728# a_472_1549# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R142 a_472_6112# m1_3338_6136# sky130_fd_pr__res_generic_m1 w=0.29 l=0.31
R143 m1_14480_5538# a_6517_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
.ends

.subckt sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2 w_415_600# a_4969_1552# a_2303_1380#
+ a_5961_1552# a_13777_1380# a_8817_1380# a_4287_1380# a_10921_1552# a_7945_1552#
+ a_12905_1552# a_7263_1380# a_12223_1380# a_9929_1552# a_9247_1380# a_2865_1380#
+ a_1993_1552# a_5841_1380# a_4849_1380# a_10801_1380# a_14135_1380# a_1311_1380#
+ a_3977_1552# a_12785_1380# a_7825_1380# a_3295_1380# a_6953_1552# a_9809_1380# a_11913_1552#
+ a_1001_1552# a_6271_1380# a_5279_1380# a_11231_1380# a_10239_1380# a_13897_1552#
+ a_8937_1552# a_8255_1380# a_1873_1380# a_13215_1380# a_3857_1380# a_2985_1552# a_11793_1380#
+ a_881_1380# a_6833_1380#
X0 a_13897_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.975 pd=6.19 as=3.775 ps=11.51 w=5 l=0.6
X1 w_415_600# a_10239_1380# a_9929_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X2 a_1993_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X3 a_8937_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X4 w_415_600# a_14135_1380# a_13897_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.72 as=2.975 ps=6.19 w=5 l=0.6
X5 w_415_600# a_3295_1380# a_2985_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X6 a_5961_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X7 w_415_600# a_2303_1380# a_1993_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X8 w_415_600# a_7263_1380# a_6953_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X9 a_4969_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X10 w_415_600# a_11231_1380# a_10921_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X11 a_12905_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X12 w_415_600# a_10239_1380# a_9929_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X13 a_8937_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X14 w_415_600# a_3295_1380# a_2985_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X15 w_415_600# a_2303_1380# a_1993_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X16 w_415_600# a_7263_1380# a_6953_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X17 a_12905_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X18 a_3977_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X19 a_7945_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X20 w_415_600# a_13215_1380# a_12905_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X21 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X22 w_415_600# a_6271_1380# a_5961_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X23 a_3977_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X24 w_415_600# a_5279_1380# a_4969_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X25 a_11913_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X26 a_7945_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X27 a_10921_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X28 w_415_600# a_13215_1380# a_12905_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X29 w_415_600# a_9247_1380# a_8937_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X30 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X31 w_415_600# a_6271_1380# a_5961_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X32 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=4.325 ps=11.73 w=5 l=0.6
X33 w_415_600# a_5279_1380# a_4969_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X34 a_11913_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X35 a_2985_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X36 a_6953_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X37 w_415_600# a_9247_1380# a_8937_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X38 a_10921_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X39 w_415_600# a_12223_1380# a_11913_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X40 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=4.325 ps=11.73 w=5 l=0.6
X41 a_9929_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X42 a_2985_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X43 w_415_600# a_4287_1380# a_3977_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X44 a_6953_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X45 w_415_600# a_8255_1380# a_7945_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X46 w_415_600# a_12223_1380# a_11913_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X47 a_13897_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.975 pd=6.19 as=3.775 ps=11.51 w=5 l=0.6
X48 a_9929_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X49 a_1993_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X50 w_415_600# a_4287_1380# a_3977_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X51 w_415_600# a_14135_1380# a_13897_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.72 as=2.975 ps=6.19 w=5 l=0.6
X52 a_5961_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
X53 w_415_600# a_11231_1380# a_10921_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X54 w_415_600# a_8255_1380# a_7945_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.775 pd=11.51 as=3.875 ps=6.55 w=5 l=0.6
X55 a_4969_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.875 pd=6.55 as=3.775 ps=11.51 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpio_pudrvr_strong_axres4v2 PU_H_N[3] PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_11913_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_8937_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_13897_1552#
+ TIE_HI_ESD sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_2985_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_4969_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_5961_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_10921_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_7945_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_12905_1552#
+ VNB sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_9929_1552# li_11868_461#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_1993_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_3977_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/w_415_600# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_6953_1552#
+ a_14575_48# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_1001_1552#
Xsky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0 sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/w_415_600#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_4969_1552# PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_5961_1552#
+ m1_14229_1478# m1_8837_1478# PU_H_N[3] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_10921_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_7945_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_12905_1552#
+ PU_H_N[3] m1_11745_1478# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_9929_1552#
+ m1_8837_1478# PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_1993_1552#
+ PU_H_N[3] PU_H_N[3] m1_10391_1478# m1_14229_1478# PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_3977_1552#
+ PU_H_N[2] PU_H_N[3] PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_6953_1552#
+ m1_10391_1478# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_11913_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_1001_1552#
+ PU_H_N[3] PU_H_N[3] m1_11745_1478# m1_10391_1478# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_13897_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_8937_1552# m1_8837_1478# PU_H_N[2]
+ m1_13667_1478# PU_H_N[3] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_2985_1552#
+ m1_11745_1478# PU_H_N[2] PU_H_N[3] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2
R0 m1_8837_1478# m2_9839_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R1 m2_14075_657# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 m1_14229_1478# m2_14532_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R3 m1_13667_1478# m2_13593_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
X0 TIE_HI_ESD a_14575_48# sky130_fd_pr__res_generic_po w=0.5 l=10.2
R4 m2_9839_n208# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 m1_10391_1478# m2_10945_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R6 m2_11422_n209# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 m1_13667_1478# m2_14075_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 m1_11745_1478# m2_12267_n279# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 m1_11745_1478# m2_12510_21# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 m2_10945_n209# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 m1_8837_1478# m2_9363_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 m1_8837_1478# m2_9605_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 m1_10391_1478# m2_11422_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 m2_9605_n209# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 m2_12510_n280# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 m2_13837_658# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 m2_14769_657# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R18 m2_11186_n208# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 m2_14286_658# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m2_14532_657# PU_H_N[3] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 m1_10391_1478# m2_11186_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 m2_13593_657# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R23 m2_12751_n280# PU_H_N[2] sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 m1_13667_1478# m2_13837_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 m1_14229_1478# m2_14769_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 m1_11745_1478# m2_12751_21# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 m2_9363_n209# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 m2_12267_n279# TIE_HI_ESD sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R29 m1_14229_1478# m2_14286_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__top_xres4v2 PAD_A_ESD_H XRES_H_N FILT_IN_H ENABLE_VDDIO TIE_WEAK_HI_H
+ ENABLE_H PULLUP_H EN_VDDIO_SIG_H TIE_LO_ESD TIE_HI_ESD DISABLE_PULLUP_H INP_SEL_H
+ VSSA VSSD AMUXBUS_B AMUXBUS_A VDDA VCCD VCCHIB VSSIO_Q VDDIO VSWITCH VSSIO PAD VDDIO_Q
Xsky130_fd_io__com_res_weak_v2_0 PULLUP_H a_5670_7125# sky130_fd_io__com_res_weak_v2
Xsky130_fd_io__com_res_weak_0 VDDIO sky130_fd_io__com_res_weak_0/RB li_7794_26629#
+ li_12154_26629# li_9658_25954# li_8568_25954# li_11000_25954# sky130_fd_io__com_res_weak
Xsky130_fd_io__xres4v2_in_buf_0 VSSD sky130_fd_io__xres4v2_in_buf_0/IN_H VDDIO_Q EN_VDDIO_SIG_H
+ sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B sky130_fd_io__xres4v2_in_buf_0/PAD ENABLE_H
+ sky130_fd_io__xres4v2_in_buf_0/IN_H_N VCCHIB ENABLE_VDDIO m1_3250_3609# EN_VDDIO_SIG_H
+ m1_1351_2970# VSSD sky130_fd_io__xres4v2_in_buf
Xsky130_fd_io__xres_inv_hysv2_0 VDDIO_Q VSSD sky130_fd_io__xres_inv_hysv2_0/OUT_H
+ m1_6377_8979# li_6043_2944# li_5552_2976# sky130_fd_io__xres_inv_hysv2
Xsky130_fd_io__gpio_buf_localesdv2_0 VSSD sky130_fd_io__xres4v2_in_buf_0/PAD sky130_fd_io__gpio_buf_localesdv2_0/OUT_VT
+ PAD VSSD VDDIO sky130_fd_io__gpio_buf_localesdv2
Xsky130_fd_io__gpio_pddrvr_strong_xres4v2_0 sky130_fd_io__gpio_pddrvr_strong_xres4v2_0/PD_H[3]
+ sky130_fd_io__gpio_pddrvr_strong_xres4v2_0/PD_H[3] sky130_fd_io__gpio_pddrvr_strong_xres4v2_0/PD_H[3]
+ VSSIO PAD PAD PAD PAD PAD PAD PAD PAD VSSIO PAD PAD PAD PAD PAD m1_915_33059# PAD
+ VDDIO sky130_fd_io__gpio_pddrvr_strong_xres4v2
Xsky130_fd_io__tk_tie_r_out_esd_0 VDDIO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd
Xsky130_fd_io__tk_tie_r_out_esd_1 VSSIO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
Xsky130_fd_io__res250only_small_0 TIE_WEAK_HI_H sky130_fd_io__com_res_weak_0/RB sky130_fd_io__res250only_small
Xsky130_fd_io__res250only_small_1 PAD PAD_A_ESD_H sky130_fd_io__res250only_small
Xsky130_fd_io__xres2v2_rcfilter_lpfv2_0 sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN
+ VDDIO_Q m1_10468_10072# m1_6377_8979# m1_10468_9216# m1_10468_4936# m1_10468_3224#
+ m1_10468_1512# m1_10468_4936# m1_10468_9216# m1_10468_3224# m1_10468_9216# m1_10468_6648#
+ m1_10468_4080# VSSD VSSD m1_10468_1512# m1_10468_7504# m1_10468_7504# m1_10468_10928#
+ m1_10468_5792# m1_10468_4080# m1_6377_8979# m1_10468_5792# m1_10468_10928# m1_10468_10072#
+ m1_10468_6648# sky130_fd_io__xres2v2_rcfilter_lpfv2
Xsky130_fd_io__gpio_pudrvr_strong_axres4v2_0 sky130_fd_io__gpio_pudrvr_strong_axres4v2_0/PU_H_N[3]
+ sky130_fd_io__gpio_pudrvr_strong_axres4v2_0/PU_H_N[3] PAD PAD PAD sky130_fd_io__gpio_pudrvr_strong_axres4v2_0/PU_H_N[3]
+ PAD PAD PAD PAD PAD PAD VSSD PAD VSSD PAD PAD VDDIO PAD VDDIO PAD sky130_fd_io__gpio_pudrvr_strong_axres4v2
X0 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 FILT_IN_H a_3226_2008# sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X2 VDDIO_Q EN_VDDIO_SIG_H sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X3 VSSD a_5525_5809# a_5551_5929# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X4 VSSD INP_SEL_H a_3226_2008# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X5 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X6 VSSD DISABLE_PULLUP_H a_5525_5809# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X7 a_5525_5809# DISABLE_PULLUP_H VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X8 a_5525_5809# DISABLE_PULLUP_H VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X9 a_3226_2008# INP_SEL_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X10 VSSD a_5556_4246# XRES_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X11 a_5551_5929# a_5525_5809# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X12 a_5556_4246# sky130_fd_io__xres_inv_hysv2_0/OUT_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X13 XRES_H_N a_5556_4246# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X14 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X15 VDDIO a_5551_5929# a_5670_7125# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.325 pd=10.53 as=0.7 ps=5.28 w=5 l=0.5
X16 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X17 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X18 VSSD a_5556_4246# XRES_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X19 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X20 XRES_H_N a_5556_4246# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X21 VDDIO_Q EN_VDDIO_SIG_H sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X22 sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X23 sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN a_3226_2008# sky130_fd_io__xres4v2_in_buf_0/IN_H VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X24 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X25 VDDIO a_5525_5809# a_5551_5929# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X26 VDDIO a_5551_5929# a_5670_7125# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X27 a_5670_7125# a_5551_5929# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X28 VDDIO DISABLE_PULLUP_H a_5525_5809# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X29 VDDIO a_5525_5809# a_5551_5929# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X30 a_3226_2008# INP_SEL_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X31 VDDIO DISABLE_PULLUP_H a_5525_5809# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X32 a_5556_4246# sky130_fd_io__xres_inv_hysv2_0/OUT_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.1855 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X33 VDDIO_Q INP_SEL_H a_3226_2008# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X34 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X35 a_5551_5929# a_5525_5809# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X36 a_5551_5929# a_5525_5809# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X37 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X38 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X39 VSSD a_5556_4246# XRES_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X40 FILT_IN_H INP_SEL_H sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X41 VSSD EN_VDDIO_SIG_H sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X42 sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X43 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X44 a_3226_2008# INP_SEL_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X45 a_5525_5809# DISABLE_PULLUP_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X46 sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN INP_SEL_H sky130_fd_io__xres4v2_in_buf_0/IN_H VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X47 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X48 VDDIO_Q INP_SEL_H a_3226_2008# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X49 VSSD a_5556_4246# XRES_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X50 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X51 a_5556_4246# sky130_fd_io__xres_inv_hysv2_0/OUT_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X52 XRES_H_N a_5556_4246# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.1855 ps=1.93 w=0.7 l=0.6
X53 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X54 sky130_fd_io__xres4v2_in_buf_0/VNORMAL_B EN_VDDIO_SIG_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X55 XRES_H_N a_5556_4246# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X56 VDDIO_Q a_5556_4246# XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X57 a_5670_7125# a_5551_5929# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.325 ps=10.53 w=5 l=0.5
X58 XRES_H_N a_5556_4246# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
.ends

.subckt sky130_ef_io__vccd_lvc_clamped_pad VDDA VCCHIB AMUXBUS_B AMUXBUS_A VCCD_PAD
+ VCCD VDDIO VSSD VSSIO VSSA VSWITCH VDDIO_Q VSSIO_Q
Xsky130_fd_io__top_power_lvc_wpad_0 VSSIO_Q VCCHIB VDDA VDDIO_Q VCCD_PAD VSSIO VSSD
+ VSSA VCCD VCCD VCCD sky130_fd_io__top_power_lvc_wpad_0/PADISOR sky130_fd_io__top_power_lvc_wpad_0/PADISOL
+ VSSA AMUXBUS_B VSSIO VDDIO VSSD VSWITCH VSSA AMUXBUS_A VCCD sky130_fd_io__top_power_lvc_wpad
.ends

.subckt sky130_fd_io__pwrdet_lshv2hv_0_pmos1 a_266_290# a_879_132# a_1191_132# w_0_0#
+ a_266_34# a_1091_34#
X0 a_879_132# a_266_290# w_0_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X1 a_266_34# a_266_290# w_0_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=2.84 as=0.42 ps=2.84 w=0.42 l=1
X2 a_266_290# a_266_34# w_0_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=2.84 as=0.42 ps=2.84 w=0.42 l=1
X3 a_1191_132# a_1091_34# w_0_0# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X4 w_0_0# a_266_290# a_879_132# w_0_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
.ends

.subckt s8_esd_res250_sub_small a_10_2# a_2142_2#
X0 a_10_2# a_2142_2# sky130_fd_pr__res_generic_po w=2 l=10.07
.ends

.subckt s8_esd_res250only_small rout pad
Xs8_esd_res250_sub_small_0 pad rout s8_esd_res250_sub_small
.ends

.subckt sky130_fd_io__pwrdet_vddd s8_esd_res250only_small_0/rout s8_esd_res250only_small_0/pad
Xs8_esd_res250only_small_0 s8_esd_res250only_small_0/rout s8_esd_res250only_small_0/pad
+ s8_esd_res250only_small
.ends

.subckt sky130_fd_io__pwrdet_vddio s8_esd_res250only_small_0/rout s8_esd_res250only_small_0/pad
Xs8_esd_res250only_small_0 s8_esd_res250only_small_0/rout s8_esd_res250only_small_0/pad
+ s8_esd_res250only_small
.ends

.subckt sky130_fd_io__pwrdet_lshv2hv_0_nmos a_65_173# a_833_141# a_1145_141# a_65_63#
+ a_1245_173# a_365_141# a_2978_173# a_2183_355# a_3086_541#
X0 a_465_173# a_365_141# a_65_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X1 a_1245_173# a_1145_141# a_1089_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X2 a_365_141# a_1145_141# a_65_63# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=1.125 pd=4.5 as=0.105 ps=1.03 w=0.75 l=0.5
X3 a_1089_173# a_833_141# a_65_63# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X4 a_1245_173# a_1145_141# a_1089_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=0.42 ps=3.28 w=3 l=0.5
X5 a_65_63# a_65_173# a_2978_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X6 a_65_173# a_365_141# a_465_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X7 a_65_63# a_2183_355# a_1145_141# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=1.125 ps=4.5 w=0.75 l=0.5
X8 a_65_63# a_833_141# a_465_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X9 a_1089_173# a_1145_141# a_1245_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X10 a_65_63# a_3086_541# a_1245_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.8
X11 a_65_63# a_1245_173# a_65_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.63 ps=3.84 w=0.42 l=1
X12 a_465_173# a_365_141# a_65_173# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=4.5 ps=9 w=3 l=0.5
X13 a_833_141# a_3086_541# a_65_63# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X14 a_1245_173# a_65_173# a_65_63# a_65_63# sky130_fd_pr__nfet_g5v0d10v5 ad=0.63 pd=3.84 as=0.0588 ps=0.7 w=0.42 l=1
.ends

.subckt sky130_fd_io__pwrdet_lshv2hv_0_pmos2 a_626_66# a_336_n32# w_100_0# a_170_66#
X0 w_100_0# a_336_n32# a_170_66# w_100_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.75 ps=3.5 w=0.75 l=0.5
X1 a_626_66# a_170_66# w_100_0# w_100_0# sky130_fd_pr__pfet_g5v0d10v5 ad=0.75 pd=3.5 as=0.105 ps=1.03 w=0.75 l=0.5
.ends

.subckt sky130_fd_io__top_pwrdetv2 in1_vddd_hv in2_vddd_hv out3_vddio_hv out1_vddio_hv
+ out2_vddio_hv out2_vddd_hv out1_vddd_hv in1_vddio_hv vddio_present_vddd_hv vddd_present_vddio_hv
+ tie_lo_esd rst_por_hv_n out3_vddd_hv in3_vddio_hv in2_vddio_hv in3_vddd_hv vssio_q
+ vccd vddd1 vssa vddio_q vddd2 vssd
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos1_0 m1_2293_2703# m1_2213_2623# m1_1977_10035#
+ vddio_q a_5004_11122# a_4058_10886# sky130_fd_io__pwrdet_lshv2hv_0_pmos1
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos1_1 m1_771_556# m1_697_476# m1_627_392# vddd1
+ a_6944_17954# a_6025_19417# sky130_fd_io__pwrdet_lshv2hv_0_pmos1
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos1_2 m1_1104_1007# m1_1032_923# m1_957_843# vddd1
+ a_6927_12695# a_6025_19417# sky130_fd_io__pwrdet_lshv2hv_0_pmos1
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos1_3 m1_4935_2408# m1_4577_2542# m1_4264_2542#
+ vddio_q a_6848_10937# a_4058_10886# sky130_fd_io__pwrdet_lshv2hv_0_pmos1
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos1_4 m1_5874_556# m1_5871_11755# m1_6663_392# vddd1
+ a_6397_12079# a_6025_19417# sky130_fd_io__pwrdet_lshv2hv_0_pmos1
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos1_5 m1_5874_2706# m1_6028_8211# m1_6663_2542#
+ vddio_q a_6848_8377# a_4058_10886# sky130_fd_io__pwrdet_lshv2hv_0_pmos1
Xsky130_fd_io__pwrdet_vddd_0 sky130_fd_io__pwrdet_vddd_0/s8_esd_res250only_small_0/rout
+ vddd2 sky130_fd_io__pwrdet_vddd
Xsky130_fd_io__pwrdet_vddio_0 sky130_fd_io__pwrdet_vddio_0/s8_esd_res250only_small_0/rout
+ vddio_q sky130_fd_io__pwrdet_vddio
Xsky130_fd_io__pwrdet_lshv2hv_0_nmos_0 m1_771_556# m1_627_392# m1_1352_1358# vssd
+ a_6944_17954# m1_1408_1468# m1_697_476# in3_vddio_hv a_6025_19417# sky130_fd_io__pwrdet_lshv2hv_0_nmos
Xsky130_fd_io__pwrdet_lshv2hv_0_nmos_1 m1_2293_2703# m1_1977_10035# m2_4976_1949#
+ vssd a_5004_11122# m1_1973_2325# m1_2213_2623# in3_vddd_hv a_4058_10886# sky130_fd_io__pwrdet_lshv2hv_0_nmos
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos2_0 m1_1408_1468# in3_vddio_hv vddio_q m1_1352_1358#
+ sky130_fd_io__pwrdet_lshv2hv_0_pmos2
Xsky130_fd_io__pwrdet_lshv2hv_0_nmos_2 m1_1104_1007# m1_957_843# m1_1520_1880# vssd
+ a_6927_12695# m1_1464_1672# m1_1032_923# in2_vddio_hv a_6025_19417# sky130_fd_io__pwrdet_lshv2hv_0_nmos
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos2_1 m1_1464_1672# in2_vddio_hv vddio_q m1_1520_1880#
+ sky130_fd_io__pwrdet_lshv2hv_0_pmos2
Xsky130_fd_io__pwrdet_lshv2hv_0_nmos_3 m1_4935_2408# m1_4264_2542# m2_5692_1949# vssd
+ a_6848_10937# m1_5621_1800# m1_4577_2542# in2_vddd_hv a_4058_10886# sky130_fd_io__pwrdet_lshv2hv_0_nmos
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos2_2 m1_1973_2325# in3_vddd_hv vddd2 m2_4976_1949#
+ sky130_fd_io__pwrdet_lshv2hv_0_pmos2
Xsky130_fd_io__pwrdet_lshv2hv_0_nmos_4 m1_5874_2706# m1_6663_2542# m2_6408_1949# vssd
+ a_6848_8377# m1_6340_1800# m1_6028_8211# in1_vddd_hv a_4058_10886# sky130_fd_io__pwrdet_lshv2hv_0_nmos
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos2_3 m1_6340_1800# in1_vddd_hv vddd2 m2_6408_1949#
+ sky130_fd_io__pwrdet_lshv2hv_0_pmos2
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos2_4 m1_5621_1800# in2_vddd_hv vddd2 m2_5692_1949#
+ sky130_fd_io__pwrdet_lshv2hv_0_pmos2
Xsky130_fd_io__pwrdet_lshv2hv_0_nmos_5 m1_5874_556# m1_6663_392# m2_3776_1949# vssd
+ a_6397_12079# m1_3708_1800# m1_5871_11755# in1_vddio_hv a_6025_19417# sky130_fd_io__pwrdet_lshv2hv_0_nmos
Xsky130_fd_io__pwrdet_lshv2hv_0_pmos2_5 m1_3708_1800# in1_vddio_hv vddio_q m2_3776_1949#
+ sky130_fd_io__pwrdet_lshv2hv_0_pmos2
X0 vssa a_2722_25404# a_3304_29317# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X1 a_3304_29317# a_2722_25404# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=10.1 ps=14.04 w=5 l=0.5
X2 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=2
X3 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X4 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X5 vddd1 a_5993_18693# vddio_present_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 a_4404_29317# rst_por_hv_n vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=2.25 ps=6 w=1.5 l=4
X7 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0 ps=0 w=1 l=4
X8 vssa vssa sky130_fd_pr__res_generic_po w=0.33 l=15.635
X9 a_3935_16143# a_2722_25404# vccd vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X10 vccd a_2722_25404# a_3935_16143# vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X11 out3_vddd_hv a_6944_18110# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X12 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0 ps=0 w=3 l=0.5
X13 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X14 a_3935_16143# a_2722_25404# vccd vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=10.5 ps=17 w=7 l=0.5
X15 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X16 vddio_present_vddd_hv a_5993_18693# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X17 out3_vddio_hv a_4985_10940# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X18 vssa a_3164_16015# a_3196_15715# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=1.5 pd=5 as=1.5 ps=5 w=1 l=8
X19 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X20 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0 ps=0 w=3 l=0.5
X21 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X22 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X23 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X24 a_5011_3767# a_4211_3735# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=4
X25 vddd1 a_6944_18110# out3_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X26 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X27 out3_vddd_hv a_6944_18110# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X28 out1_vddd_hv a_6378_12177# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X29 vssd a_6927_12695# a_6817_12995# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X30 vssd a_6848_9735# out2_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X31 vssa a_4211_3735# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X32 vssa a_2722_25404# a_3935_14683# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=4.5 ps=9 w=3 l=8
X33 vddd1 a_6378_12177# out1_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X34 a_3304_29317# a_3164_16015# a_4404_29317# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=2.25 pd=6 as=0.21 ps=1.78 w=1.5 l=4
X35 out2_vddd_hv a_6817_12995# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X36 out2_vddd_hv a_6817_12995# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X37 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X38 a_3634_17232# a_3196_15715# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X39 out3_vddd_hv a_6944_18110# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X40 out2_vddio_hv a_6848_9735# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X41 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X42 out1_vddd_hv a_6378_12177# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X43 vddio_q a_3144_11068# a_4058_10886# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.56 as=0.21 ps=1.78 w=1.5 l=0.5
X44 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X45 out1_vddio_hv a_6848_9111# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X46 vssd a_3634_17232# a_6025_19417# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X47 vssd a_6944_17954# a_6944_18110# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X48 vddd_present_vddio_hv a_3122_10886# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X49 a_3144_11068# a_5011_3767# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=2
X50 a_4058_10886# a_3144_11068# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X51 vssd a_6817_12995# out2_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X52 out1_vddio_hv a_6848_9111# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X53 out3_vddio_hv a_4985_10940# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X54 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X55 vddio_q a_3122_10886# vddd_present_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X56 vddd1 a_6927_12695# a_6817_12995# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X57 out2_vddio_hv a_6848_9735# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X58 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0 ps=0 w=1 l=8
X59 a_6025_19417# a_3634_17232# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X60 vddd1 a_6397_12079# a_6378_12177# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X61 a_4404_29317# a_3164_16015# a_3304_29317# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=2.25 ps=6 w=1.5 l=4
X62 vddio_present_vddd_hv a_5993_18693# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X63 vssd a_5993_18693# vddio_present_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X64 vddio_q a_5004_11122# a_4985_10940# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X65 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X66 vddio_q a_3122_10886# vddd_present_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X67 a_3208_7281# a_3039_3259# a_3139_3291# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=4.5 ps=9 w=3 l=8
X68 vddd1 a_3634_17232# a_6025_19417# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X69 tie_lo_esd vssd sky130_fd_pr__res_generic_po w=0.5 l=10.2
X70 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.5
X71 vssa a_3935_16143# a_3164_16015# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7.5 pd=13 as=0.7 ps=5.28 w=5 l=0.5
X72 a_2352_39489# a_9590_39549# sky130_fd_pr__res_generic_po w=0.33 l=1.95k
X73 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0 ps=0 w=3 l=0.5
X74 out3_vddd_hv a_6944_18110# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X75 vssd a_4985_10940# out3_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X76 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0 ps=0 w=3 l=0.5
X77 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0 ps=0 w=3 l=0.5
X78 a_5011_3767# a_4211_3735# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=4
X79 vddd1 a_3164_16015# a_3196_15715# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=1.5 pd=5 as=0.14 ps=1.28 w=1 l=8
X80 vddio_present_vddd_hv a_5993_18693# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X81 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0 ps=0 w=3 l=0.5
X82 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0 ps=0 w=3 l=0.5
X83 vddd1 a_6817_12995# out2_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X84 a_3139_3291# a_3039_3259# a_552_39489# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X85 a_6848_9111# a_6848_8377# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X86 out2_vddd_hv a_6817_12995# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X87 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X88 vccd a_2722_25404# a_3935_16143# vccd sky130_fd_pr__pfet_g5v0d10v5 ad=10.5 pd=17 as=0.98 ps=7.28 w=7 l=0.5
X89 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X90 vddd1 a_6944_18110# out3_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X91 vddd1 a_6944_18110# out3_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X92 vssd a_6944_18110# out3_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X93 vddd1 a_6378_12177# out1_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X94 vssd a_6397_12079# a_6378_12177# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X95 vssd a_6848_9111# out1_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X96 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X97 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X98 out3_vddio_hv a_4985_10940# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X99 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X100 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X101 vddio_q a_6848_9111# out1_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X102 vddio_q a_4985_10940# out3_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X103 out2_vddio_hv a_6848_9735# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X104 vddd1 a_6817_12995# out2_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X105 vddd1 a_3196_15715# a_3634_17232# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X106 vssa a_3196_15715# a_3634_17232# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0.105 ps=1.03 w=0.75 l=0.5
X107 vssa a_3039_3259# a_3938_5381# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=4.5 ps=9 w=3 l=8
X108 vssd a_6378_12177# out1_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X109 vddd1 a_6944_17954# a_6944_18110# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X110 vddio_q a_6848_9735# out2_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X111 out1_vddd_hv a_6378_12177# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X112 out1_vddd_hv a_6378_12177# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X113 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X114 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X115 vssd a_3144_11068# a_4058_10886# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0.105 ps=1.03 w=0.75 l=0.5
X116 a_6025_19417# a_3634_17232# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X117 out2_vddd_hv a_6817_12995# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X118 a_4058_10886# a_3144_11068# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X119 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X120 vssa a_4211_3735# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X121 a_3634_17232# a_3196_15715# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X122 vddio_q a_6848_9111# out1_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X123 vddio_q a_4211_3735# a_5011_3767# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=4
X124 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X125 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X126 vssa a_4211_3735# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X127 vddd2 vddd2 vssd sky130_fd_pr__res_generic_nd__hv w=0.3 l=68.84
X128 vssa a_4211_3735# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X129 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0 ps=0 w=0.75 l=0.5
X130 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0 ps=0 w=1.5 l=0.5
X131 vddio_q a_5011_3767# a_3144_11068# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=2
X132 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0 ps=0 w=0.75 l=0.5
X133 vssd a_6378_12177# out1_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X134 vssa a_4211_3735# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X135 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0 ps=0 w=0.75 l=0.5
X136 a_3304_29317# rst_por_hv_n vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=1.5 pd=5 as=1.5 ps=5 w=1 l=1
X137 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X138 out1_vddd_hv a_6378_12177# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X139 vssd a_3144_11068# a_4058_10886# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X140 a_3164_16015# a_3935_16143# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X141 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0 ps=0 w=1.5 l=0.5
X142 vssd a_3122_10886# vddd_present_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X143 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0 ps=0 w=3 l=0.5
X144 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0 ps=0 w=3 l=0.5
X145 vddd1 a_3634_17232# a_5993_18693# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.42 ps=3.56 w=1.5 l=0.5
X146 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0 ps=0 w=1.5 l=0.5
X147 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X148 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0 ps=0 w=3 l=0.5
X149 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0 ps=0 w=0.75 l=0.5
X150 a_552_39489# a_3039_3259# a_3139_3291# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X151 out3_vddd_hv a_6944_18110# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X152 a_3139_3291# a_3039_3259# a_552_39489# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=10.395 ps=16.97 w=7 l=0.5
X153 out2_vddio_hv a_6848_9735# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X154 vddd1 a_6378_12177# out1_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X155 out2_vddio_hv a_6848_9735# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X156 vssd a_3634_17232# a_6025_19417# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=2.06 as=0.105 ps=1.03 w=0.75 l=0.5
X157 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X158 out3_vddio_hv a_4985_10940# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X159 vssd a_6848_9735# out2_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X160 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X161 out1_vddio_hv a_6848_9111# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X162 out1_vddio_hv a_6848_9111# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X163 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.5
X164 a_3164_16015# a_3935_16143# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X165 a_9590_39549# vddio_q vssd sky130_fd_pr__res_generic_nd__hv w=0.3 l=1.33932k
X166 a_3304_29317# a_2722_25404# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X167 vddio_q a_6848_9735# out2_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X168 a_3208_7281# a_3039_3259# a_3938_5381# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=4.5 ps=9 w=3 l=8
X169 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.56 as=0 ps=0 w=10 l=2
X170 vssa a_3935_16143# a_3164_16015# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X171 out1_vddd_hv a_6378_12177# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X172 out2_vddio_hv a_6848_9735# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X173 a_4058_10886# a_3144_11068# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X174 vssa vssa vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0 ps=0 w=1 l=4
X175 vddd1 a_6378_12177# out1_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X176 vddio_q a_4985_10940# out3_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X177 out2_vddd_hv a_6817_12995# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X178 out2_vddd_hv a_6817_12995# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X179 vddio_q a_6848_8377# a_6848_9111# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X180 vssa a_3304_29317# a_3164_16015# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=2.25 pd=6 as=0.21 ps=1.78 w=1.5 l=4
X181 a_3935_16143# a_2722_25404# vccd vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X182 a_3634_17232# a_3196_15715# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21 ps=2.06 w=0.75 l=0.5
X183 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X184 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X185 vccd a_2722_25404# a_3935_16143# vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X186 vddd1 a_3634_17232# a_6025_19417# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.56 as=0.21 ps=1.78 w=1.5 l=0.5
X187 out3_vddd_hv a_6944_18110# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X188 vddio_q a_3144_11068# a_4058_10886# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X189 vddd_present_vddio_hv a_3122_10886# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X190 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X191 vssd a_5993_18693# vddio_present_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X192 out1_vddio_hv a_6848_9111# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X193 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X194 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X195 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X196 vssd a_6817_12995# out2_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X197 vddio_present_vddd_hv a_5993_18693# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X198 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X199 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X200 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.56 as=0 ps=0 w=1.5 l=0.5
X201 vssd a_3122_10886# vddd_present_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X202 a_6025_19417# a_3634_17232# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X203 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0 ps=0 w=1.5 l=0.5
X204 vddd_present_vddio_hv a_3122_10886# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X205 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0 ps=0 w=3 l=0.5
X206 vddd1 a_3164_16015# a_3304_29317# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.63 pd=3.84 as=0.63 ps=3.84 w=0.42 l=20
X207 vssd a_3634_17232# a_5993_18693# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21 ps=2.06 w=0.75 l=0.5
X208 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X209 a_3164_16015# a_3304_29317# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=2.25 ps=6 w=1.5 l=4
X210 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0 ps=0 w=3 l=0.5
X211 vssd a_6944_18110# out3_vddd_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X212 a_552_39489# a_3039_3259# a_3139_3291# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=10.5 pd=17 as=0.98 ps=7.28 w=7 l=0.5
X213 vssd a_5004_11122# a_4985_10940# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X214 a_5835_15413# a_2722_25404# a_3935_16143# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=4.5 ps=9 w=3 l=8
X215 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0 ps=0 w=3 l=0.5
X216 a_3935_16143# a_2722_25404# vccd vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X217 vddd1 a_5993_18693# vddio_present_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X218 vddio_q a_4985_10940# out3_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X219 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X220 vssd a_4985_10940# out3_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X221 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X222 vddd1 vddd1 vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.56 as=0 ps=0 w=1.5 l=0.5
X223 vddio_q a_6848_9111# out1_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X224 a_5835_15413# a_2722_25404# a_3935_14683# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=4.5 pd=9 as=4.5 ps=9 w=3 l=8
X225 a_4211_3735# a_3139_3291# a_3967_4161# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=1.5 pd=5 as=1.5 ps=5 w=1 l=8
X226 out3_vddio_hv a_4985_10940# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X227 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X228 a_3039_3259# sky130_fd_io__pwrdet_vddd_0/s8_esd_res250only_small_0/rout vssd sky130_fd_pr__res_generic_nd__hv w=0.3 l=68.84
X229 vddio_q a_6848_9735# out2_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X230 vddio_q a_6848_9735# out2_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X231 out3_vddio_hv a_4985_10940# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X232 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X233 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0 ps=0 w=1.5 l=0.5
X234 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X235 vddio_q a_4985_10940# out3_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X236 vssa a_5011_3767# a_3144_11068# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=2
X237 vddd1 a_3304_29317# a_3164_16015# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.63 pd=3.84 as=0.63 ps=3.84 w=0.42 l=20
X238 vssa a_2722_25404# a_3304_29317# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X239 vddd1 a_6817_12995# out2_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X240 out1_vddio_hv a_6848_9111# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X241 vddd_present_vddio_hv a_3122_10886# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X242 vssa a_3196_15715# a_3634_17232# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X243 vssd a_3144_11068# a_3122_10886# vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.21 ps=2.06 w=0.75 l=0.5
X244 a_3196_15715# a_3164_16015# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=1.5 ps=5 w=1 l=8
X245 vddd1 a_6944_18110# out3_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X246 a_6848_9735# a_6848_10937# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.19875 ps=2.03 w=0.75 l=0.5
X247 vssd a_6848_9111# out1_vddio_hv vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X248 a_4211_3735# a_3139_3291# vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=7.7 pd=16.2 as=7.7 ps=16.2 w=7 l=0.5
X249 vssa rst_por_hv_n a_4404_29317# vssa sky130_fd_pr__nfet_g5v0d10v5 ad=2.25 pd=6 as=0.21 ps=1.78 w=1.5 l=4
X250 vddio_q a_6848_9111# out1_vddio_hv vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X251 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X252 vccd a_2722_25404# a_3935_16143# vccd sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X253 vddd1 a_6817_12995# out2_vddd_hv vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X254 a_552_39489# a_2352_39489# vssd sky130_fd_pr__res_generic_nd__hv w=0.3 l=3.14938k
X255 vddd1 a_3196_15715# a_3634_17232# vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X256 vddio_q a_6848_10937# a_6848_9735# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X257 vssd vssd vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X258 a_6025_19417# a_3634_17232# vssd vssd sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X259 a_4058_10886# a_3144_11068# vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X260 vddio_q a_3144_11068# a_3122_10886# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.42 ps=3.56 w=1.5 l=0.5
X261 vssa a_2722_25404# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X262 vssa a_3039_3259# vssa vssa sky130_fd_pr__nfet_05v0_nvt ad=1.4 pd=10.28 as=0 ps=0 w=10 l=2
X263 a_2722_25404# sky130_fd_io__pwrdet_vddio_0/s8_esd_res250only_small_0/rout vssd sky130_fd_pr__res_generic_nd__hv w=0.3 l=277.39001
X264 vddio_q vddio_q vddio_q vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0 ps=0 w=1.5 l=0.5
X265 a_3634_17232# a_3196_15715# vddd1 vddd1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X266 vddio_q a_3139_3291# a_3967_4161# vddio_q sky130_fd_pr__pfet_g5v0d10v5 ad=1.5 pd=5 as=1.5 ps=5 w=1 l=8
.ends

.subckt sky130_ef_io__vssd_lvc_clamped_pad VDDA VSSD_PAD VCCD VSWITCH VDDIO AMUXBUS_A
+ AMUXBUS_B VDDIO_Q VSSD VSSIO VSSIO_Q VCCHIB VSSA
Xsky130_fd_io__top_ground_lvc_wpad_1 sky130_fd_io__top_ground_lvc_wpad_1/PADISOR sky130_fd_io__top_ground_lvc_wpad_1/PADISOL
+ VSSIO_Q VCCHIB VDDA VDDIO_Q VSSD_PAD VSSIO VSSD VSSA VCCD VCCD VSSD VSSA AMUXBUS_B
+ VSSIO VDDIO VSSD VSWITCH VSSA AMUXBUS_A VCCD sky130_fd_io__top_ground_lvc_wpad
.ends

.subckt panamax vccd0_0 select resetb gpio8_0 gpio8_1 gpio8_2 gpio8_3 vssio_8 vssd0_0
+ xi0 xo0 xi1 xo1 vddio_9 vccd0_1 gpio8_4 gpio8_5 gpio8_6 gpio8_7 vssio_9 vssa3_0
+ vdda3_0 vssd0_1 sio0 sio1 vddio_0 gpio0_0 gpio0_1 gpio0_2 gpio0_3 vssd1_0 vssio_0
+ gpio0_4 gpio0_5 gpio0_6 gpio0_7 vddio_1 vdda1_0 vssa1_0 gpio1_0 gpio1_1 gpio1_2
+ gpio1_3 vccd1_0 vssio_1 gpio1_4 gpio1_5 gpio1_6 gpio1_7 vddio_2 vdda1_1 vssa1_1
+ vssd1_1 gpio2_0 gpio2_1 gpio2_2 gpio2_3 vssio_2 gpio2_4 gpio2_5 gpio2_6 gpio2_7
+ vccd1_1 vddio_3 vccd2_0 gpio4_7 gpio4_6 gpio4_5 gpio4_4 vssio_4 vssd2_0 gpio4_3
+ gpio4_2 gpio4_1 gpio4_0 vssa0_0 analog_1 analog_0 vdda0_0 vddio_4 gpio3_7 gpio3_6
+ gpio3_5 gpio3_4 vccd1_2 vssio_3 gpio3_3 gpio3_2 gpio3_1 gpio3_0 vssd1_2 vddio_8
+ gpio7_7 gpio7_6 gpio7_5 gpio7_4 vccd2_2 vssio_7 gpio7_3 gpio7_2 gpio7_1 gpio7_0
+ vddio_7 vdda2_1 vssa2_1 gpio6_7 gpio6_6 gpio6_5 gpio6_4 vssd2_2 vssio_6 gpio6_3
+ gpio6_2 gpio6_1 gpio6_0 vddio_6 vdda2_0 vssa2_0 vccd2_1 gpio5_7 gpio5_6 gpio5_5
+ gpio5_4 vssio_5 gpio5_3 gpio5_2 gpio5_1 gpio5_0 vssd2_1 vddio_5 vccd0 vssio vssd0
+ vddio vssa3 vdda3 vssd1[0] vccd1[0] vdda1 vssa1 vccd1[1] vssd1[1] vssd1[2] vccd1[2]
+ vccd1[3] vssd1[3] vssd1[4] vccd1[4] vccd1[5] vssd1[5] vdda0 vssa0 vssd2[0] vccd2[0]
+ vccd2[1] vssd2[1] vssd2[2] vccd2[2] vccd2[3] vssd2[3] vssa2 vdda2 vssd2[4] vccd2[4]
+ vccd2[5] vssd2[5] select_tie_lo_esd select_in select_tie_hi_esd select_enable_vddio
+ select_slow select_pad_a_esd_0_h select_pad_a_esd_1_h select_pad_a_noesd_h select_analog_en
+ select_analog_pol select_inp_dis select_enable_inp_h select_enable_h select_hld_h_n
+ select_analog_sel select_dm[2] select_dm[1] select_dm[0] select_hld_ovr select_out
+ select_enable_vswitch_h select_enable_vdda_h select_vtrip_sel select_ib_mode_sel
+ select_oe_n select_in_h select_zero select_one resetb_tie_weak_hi_h resetb_disable_pullup_h
+ resetb_tie_hi_esd resetb_xres_h_n resetb_tie_lo_esd resetb_inp_sel_h resetb_en_vddio_sig_h
+ resetb_filt_in_h resetb_pad_a_esd_h resetb_pullup_h resetb_enable_h resetb_enable_vddio
+ gpio8_0_tie_lo_esd gpio8_0_in gpio8_0_tie_hi_esd gpio8_0_enable_vddio gpio8_0_slow
+ gpio8_0_pad_a_esd_0_h gpio8_0_pad_a_esd_1_h gpio8_0_pad_a_noesd_h gpio8_0_analog_en
+ gpio8_0_analog_pol gpio8_0_inp_dis gpio8_0_enable_inp_h gpio8_0_enable_h gpio8_0_hld_h_n
+ gpio8_0_analog_sel gpio8_0_dm[2] gpio8_0_dm[1] gpio8_0_dm[0] gpio8_0_hld_ovr gpio8_0_out
+ gpio8_0_enable_vswitch_h gpio8_0_enable_vdda_h gpio8_0_vtrip_sel gpio8_0_ib_mode_sel
+ gpio8_0_oe_n gpio8_0_in_h gpio8_0_zero gpio8_0_one gpio8_1_tie_lo_esd gpio8_1_in
+ gpio8_1_tie_hi_esd gpio8_1_enable_vddio gpio8_1_slow gpio8_1_pad_a_esd_0_h gpio8_1_pad_a_esd_1_h
+ gpio8_1_pad_a_noesd_h gpio8_1_analog_en gpio8_1_analog_pol gpio8_1_inp_dis gpio8_1_enable_inp_h
+ gpio8_1_enable_h gpio8_1_hld_h_n gpio8_1_analog_sel gpio8_1_dm[2] gpio8_1_dm[1]
+ gpio8_1_dm[0] gpio8_1_hld_ovr gpio8_1_out gpio8_1_enable_vswitch_h gpio8_1_enable_vdda_h
+ gpio8_1_vtrip_sel gpio8_1_ib_mode_sel gpio8_1_oe_n gpio8_1_in_h gpio8_1_zero gpio8_1_one
+ gpio8_2_tie_lo_esd gpio8_2_in gpio8_2_tie_hi_esd gpio8_2_enable_vddio gpio8_2_slow
+ gpio8_2_pad_a_esd_0_h gpio8_2_pad_a_esd_1_h gpio8_2_pad_a_noesd_h gpio8_2_analog_en
+ gpio8_2_analog_pol gpio8_2_inp_dis gpio8_2_enable_inp_h gpio8_2_enable_h gpio8_2_hld_h_n
+ gpio8_2_analog_sel gpio8_2_dm[2] gpio8_2_dm[1] gpio8_2_dm[0] gpio8_2_hld_ovr gpio8_2_out
+ gpio8_2_enable_vswitch_h gpio8_2_enable_vdda_h gpio8_2_vtrip_sel gpio8_2_ib_mode_sel
+ gpio8_2_oe_n gpio8_2_in_h gpio8_2_zero gpio8_2_one gpio8_3_tie_lo_esd gpio8_3_in
+ gpio8_3_tie_hi_esd gpio8_3_enable_vddio gpio8_3_slow gpio8_3_pad_a_esd_0_h gpio8_3_pad_a_esd_1_h
+ gpio8_3_pad_a_noesd_h gpio8_3_analog_en gpio8_3_analog_pol gpio8_3_inp_dis gpio8_3_enable_inp_h
+ gpio8_3_enable_h gpio8_3_hld_h_n gpio8_3_analog_sel gpio8_3_dm[2] gpio8_3_dm[1]
+ gpio8_3_dm[0] gpio8_3_hld_ovr gpio8_3_out gpio8_3_enable_vswitch_h gpio8_3_enable_vdda_h
+ gpio8_3_vtrip_sel gpio8_3_ib_mode_sel gpio8_3_oe_n gpio8_3_in_h gpio8_3_zero gpio8_3_one
+ xi0_core xo0_core xi1_core xo1_core gpio8_4_tie_lo_esd gpio8_4_in gpio8_4_tie_hi_esd
+ gpio8_4_enable_vddio gpio8_4_slow gpio8_4_pad_a_esd_0_h gpio8_4_pad_a_esd_1_h gpio8_4_pad_a_noesd_h
+ gpio8_4_analog_en gpio8_4_analog_pol gpio8_4_inp_dis gpio8_4_enable_inp_h gpio8_4_enable_h
+ gpio8_4_hld_h_n gpio8_4_analog_sel gpio8_4_dm[2] gpio8_4_dm[1] gpio8_4_dm[0] gpio8_4_hld_ovr
+ gpio8_4_out gpio8_4_enable_vswitch_h gpio8_4_enable_vdda_h gpio8_4_vtrip_sel gpio8_4_ib_mode_sel
+ gpio8_4_oe_n gpio8_4_in_h gpio8_4_zero gpio8_4_one gpio8_5_tie_lo_esd gpio8_5_in
+ gpio8_5_tie_hi_esd gpio8_5_enable_vddio gpio8_5_slow gpio8_5_pad_a_esd_0_h gpio8_5_pad_a_esd_1_h
+ gpio8_5_pad_a_noesd_h gpio8_5_analog_en gpio8_5_analog_pol gpio8_5_inp_dis gpio8_5_enable_inp_h
+ gpio8_5_enable_h gpio8_5_hld_h_n gpio8_5_analog_sel gpio8_5_dm[2] gpio8_5_dm[1]
+ gpio8_5_dm[0] gpio8_5_hld_ovr gpio8_5_out gpio8_5_enable_vswitch_h gpio8_5_enable_vdda_h
+ gpio8_5_vtrip_sel gpio8_5_ib_mode_sel gpio8_5_oe_n gpio8_5_in_h gpio8_5_zero gpio8_5_one
+ gpio8_6_tie_lo_esd gpio8_6_in gpio8_6_tie_hi_esd gpio8_6_enable_vddio gpio8_6_slow
+ gpio8_6_pad_a_esd_0_h gpio8_6_pad_a_esd_1_h gpio8_6_pad_a_noesd_h gpio8_6_analog_en
+ gpio8_6_analog_pol gpio8_6_inp_dis gpio8_6_enable_inp_h gpio8_6_enable_h gpio8_6_hld_h_n
+ gpio8_6_analog_sel gpio8_6_dm[2] gpio8_6_dm[1] gpio8_6_dm[0] gpio8_6_hld_ovr gpio8_6_out
+ gpio8_6_enable_vswitch_h gpio8_6_enable_vdda_h gpio8_6_vtrip_sel gpio8_6_ib_mode_sel
+ gpio8_6_oe_n gpio8_6_in_h gpio8_6_zero gpio8_6_one gpio8_7_tie_lo_esd gpio8_7_in
+ gpio8_7_tie_hi_esd gpio8_7_enable_vddio gpio8_7_slow gpio8_7_pad_a_esd_0_h gpio8_7_pad_a_esd_1_h
+ gpio8_7_pad_a_noesd_h gpio8_7_analog_en gpio8_7_analog_pol gpio8_7_inp_dis gpio8_7_enable_inp_h
+ gpio8_7_enable_h gpio8_7_hld_h_n gpio8_7_analog_sel gpio8_7_dm[2] gpio8_7_dm[1]
+ gpio8_7_dm[0] gpio8_7_hld_ovr gpio8_7_out gpio8_7_enable_vswitch_h gpio8_7_enable_vdda_h
+ gpio8_7_vtrip_sel gpio8_7_ib_mode_sel gpio8_7_oe_n gpio8_7_in_h gpio8_7_zero gpio8_7_one
+ pwrdet_out2_vddio_hv pwrdet_out1_vddd_hv pwrdet_in1_vddio_hv pwrdet_in2_vddd_hv
+ pwrdet_in1_vddd_hv pwrdet_out1_vddio_hv pwrdet_out2_vddd_hv pwrdet_out3_vddd_hv
+ pwrdet_vddio_present_vddd_hv pwrdet_out3_vddio_hv pwrdet_tie_lo_esd pwrdet_in3_vddd_hv
+ pwrdet_vddd_present_vddio_hv pwrdet_in2_vddio_hv pwrdet_in3_vddio_hv pwrdet_rst_por_hv_n
+ sio_vinref_dft sio_voutref_dft sio_vref_sel[1] sio_vref_sel[0] sio_enable_vdda_h
+ sio_dft_refgen sio_voh_sel[2] sio_voh_sel[1] sio_voh_sel[0] amuxbus_a_n amuxbus_b_n
+ sio_amuxbus_b sio_amuxbus_a sio_vreg_en_refgen sio_ibuf_sel_refgen sio_vohref sio_hld_h_n_refgen
+ sio_vtrip_sel_refgen sio_pad_a_esd_0_h[1] sio_pad_a_noesd_h[1] sio_inp_dis[1] sio_tie_lo_esd[1]
+ sio_out[1] sio_vtrip_sel[1] sio_ibuf_sel[1] sio_hld_h_n[1] sio_hld_ovr[1] sio_in[1]
+ sio_in_h[1] sio_oe_n[1] sio_slow[1] sio_vreg_en[1] sio_enable_h sio_dm1[2] sio_dm1[1]
+ sio_dm1[0] sio_pad_a_esd_1_h[1] sio_pad_a_esd_1_h[0] sio_dm0[0] sio_dm0[1] sio_dm0[2]
+ sio_vreg_en[0] sio_slow[0] sio_oe_n[0] sio_in_h[0] sio_in[0] sio_hld_ovr[0] sio_hld_h_n[0]
+ sio_ibuf_sel[0] sio_vtrip_sel[0] sio_out[0] sio_tie_lo_esd[0] sio_inp_dis[0] sio_pad_a_noesd_h[0]
+ sio_pad_a_esd_0_h[0] muxsplit_se_hld_vdda_h_n muxsplit_se_enable_vdda_h muxsplit_se_switch_aa_sl
+ muxsplit_se_switch_aa_s0 muxsplit_se_switch_bb_s0 muxsplit_se_switch_bb_sl muxsplit_se_switch_bb_sr
+ muxsplit_se_switch_aa_sr gpio0_0_tie_lo_esd gpio0_0_in gpio0_0_tie_hi_esd gpio0_0_enable_vddio
+ gpio0_0_slow gpio0_0_pad_a_esd_0_h gpio0_0_pad_a_esd_1_h gpio0_0_pad_a_noesd_h gpio0_0_analog_en
+ gpio0_0_analog_pol gpio0_0_inp_dis gpio0_0_enable_inp_h gpio0_0_enable_h gpio0_0_hld_h_n
+ gpio0_0_analog_sel gpio0_0_dm[2] gpio0_0_dm[1] gpio0_0_dm[0] gpio0_0_hld_ovr gpio0_0_out
+ gpio0_0_enable_vswitch_h gpio0_0_enable_vdda_h gpio0_0_vtrip_sel gpio0_0_ib_mode_sel
+ gpio0_0_oe_n gpio0_0_in_h gpio0_0_zero gpio0_0_one gpio0_1_tie_lo_esd gpio0_1_in
+ gpio0_1_tie_hi_esd gpio0_1_enable_vddio gpio0_1_slow gpio0_1_pad_a_esd_0_h gpio0_1_pad_a_esd_1_h
+ gpio0_1_pad_a_noesd_h gpio0_1_analog_en gpio0_1_analog_pol gpio0_1_inp_dis gpio0_1_enable_inp_h
+ gpio0_1_enable_h gpio0_1_hld_h_n gpio0_1_analog_sel gpio0_1_dm[2] gpio0_1_dm[1]
+ gpio0_1_dm[0] gpio0_1_hld_ovr gpio0_1_out gpio0_1_enable_vswitch_h gpio0_1_enable_vdda_h
+ gpio0_1_vtrip_sel gpio0_1_ib_mode_sel gpio0_1_oe_n gpio0_1_in_h gpio0_1_zero gpio0_1_one
+ gpio0_2_tie_lo_esd gpio0_2_in gpio0_2_tie_hi_esd gpio0_2_enable_vddio gpio0_2_slow
+ gpio0_2_pad_a_esd_0_h gpio0_2_pad_a_esd_1_h gpio0_2_pad_a_noesd_h gpio0_2_analog_en
+ gpio0_2_analog_pol gpio0_2_inp_dis gpio0_2_enable_inp_h gpio0_2_enable_h gpio0_2_hld_h_n
+ gpio0_2_analog_sel gpio0_2_dm[2] gpio0_2_dm[1] gpio0_2_dm[0] gpio0_2_hld_ovr gpio0_2_out
+ gpio0_2_enable_vswitch_h gpio0_2_enable_vdda_h gpio0_2_vtrip_sel gpio0_2_ib_mode_sel
+ gpio0_2_oe_n gpio0_2_in_h gpio0_2_zero gpio0_2_one gpio0_3_tie_lo_esd gpio0_3_in
+ gpio0_3_tie_hi_esd gpio0_3_enable_vddio gpio0_3_slow gpio0_3_pad_a_esd_0_h gpio0_3_pad_a_esd_1_h
+ gpio0_3_pad_a_noesd_h gpio0_3_analog_en gpio0_3_analog_pol gpio0_3_inp_dis gpio0_3_enable_inp_h
+ gpio0_3_enable_h gpio0_3_hld_h_n gpio0_3_analog_sel gpio0_3_dm[2] gpio0_3_dm[1]
+ gpio0_3_dm[0] gpio0_3_hld_ovr gpio0_3_out gpio0_3_enable_vswitch_h gpio0_3_enable_vdda_h
+ gpio0_3_vtrip_sel gpio0_3_ib_mode_sel gpio0_3_oe_n gpio0_3_in_h gpio0_3_zero gpio0_3_one
+ gpio0_4_tie_lo_esd gpio0_4_in gpio0_4_tie_hi_esd gpio0_4_enable_vddio gpio0_4_slow
+ gpio0_4_pad_a_esd_0_h gpio0_4_pad_a_esd_1_h gpio0_4_pad_a_noesd_h gpio0_4_analog_en
+ gpio0_4_analog_pol gpio0_4_inp_dis gpio0_4_enable_inp_h gpio0_4_enable_h gpio0_4_hld_h_n
+ gpio0_4_analog_sel gpio0_4_dm[2] gpio0_4_dm[1] gpio0_4_dm[0] gpio0_4_hld_ovr gpio0_4_out
+ gpio0_4_enable_vswitch_h gpio0_4_enable_vdda_h gpio0_4_vtrip_sel gpio0_4_ib_mode_sel
+ gpio0_4_oe_n gpio0_4_in_h gpio0_4_zero gpio0_4_one gpio0_5_tie_lo_esd gpio0_5_in
+ gpio0_5_tie_hi_esd gpio0_5_enable_vddio gpio0_5_slow gpio0_5_pad_a_esd_0_h gpio0_5_pad_a_esd_1_h
+ gpio0_5_pad_a_noesd_h gpio0_5_analog_en gpio0_5_analog_pol gpio0_5_inp_dis gpio0_5_enable_inp_h
+ gpio0_5_enable_h gpio0_5_hld_h_n gpio0_5_analog_sel gpio0_5_dm[2] gpio0_5_dm[1]
+ gpio0_5_dm[0] gpio0_5_hld_ovr gpio0_5_out gpio0_5_enable_vswitch_h gpio0_5_enable_vdda_h
+ gpio0_5_vtrip_sel gpio0_5_ib_mode_sel gpio0_5_oe_n gpio0_5_in_h gpio0_5_zero gpio0_5_one
+ gpio0_6_tie_lo_esd gpio0_6_in gpio0_6_tie_hi_esd gpio0_6_enable_vddio gpio0_6_slow
+ gpio0_6_pad_a_esd_0_h gpio0_6_pad_a_esd_1_h gpio0_6_pad_a_noesd_h gpio0_6_analog_en
+ gpio0_6_analog_pol gpio0_6_inp_dis gpio0_6_enable_inp_h gpio0_6_enable_h gpio0_6_hld_h_n
+ gpio0_6_analog_sel gpio0_6_dm[2] gpio0_6_dm[1] gpio0_6_dm[0] gpio0_6_hld_ovr gpio0_6_out
+ gpio0_6_enable_vswitch_h gpio0_6_enable_vdda_h gpio0_6_vtrip_sel gpio0_6_ib_mode_sel
+ gpio0_6_oe_n gpio0_6_in_h gpio0_6_zero gpio0_6_one gpio0_7_tie_lo_esd gpio0_7_in
+ gpio0_7_tie_hi_esd gpio0_7_enable_vddio gpio0_7_slow gpio0_7_pad_a_esd_0_h gpio0_7_pad_a_esd_1_h
+ gpio0_7_pad_a_noesd_h gpio0_7_analog_en gpio0_7_analog_pol gpio0_7_inp_dis gpio0_7_enable_inp_h
+ gpio0_7_enable_h gpio0_7_hld_h_n gpio0_7_analog_sel gpio0_7_dm[2] gpio0_7_dm[1]
+ gpio0_7_dm[0] gpio0_7_hld_ovr gpio0_7_out gpio0_7_enable_vswitch_h gpio0_7_enable_vdda_h
+ gpio0_7_vtrip_sel gpio0_7_ib_mode_sel gpio0_7_oe_n gpio0_7_in_h gpio0_7_zero gpio0_7_one
+ gpio1_0_tie_hi_esd gpio1_0_dm[2] gpio1_0_dm[1] gpio1_0_dm[0] gpio1_0_slow gpio1_0_oe_n
+ gpio1_0_tie_lo_esd gpio1_0_inp_dis gpio1_0_enable_vddio gpio1_0_vtrip_sel gpio1_0_ib_mode_sel[1]
+ gpio1_0_ib_mode_sel[0] gpio1_0_out gpio1_0_slew_ctl[1] gpio1_0_slew_ctl[0] gpio1_0_analog_pol
+ gpio1_0_analog_sel gpio1_0_hys_trim gpio1_0_hld_ovr gpio1_0_in_h gpio1_0_enable_h
+ gpio1_0_in gpio1_0_hld_h_n gpio1_0_enable_vdda_h gpio1_0_analog_en gpio1_0_enable_inp_h
+ gpio1_0_enable_vswitch_h gpio1_0_pad_a_noesd_h gpio1_0_pad_a_esd_0_h gpio1_0_pad_a_esd_1_h
+ gpio1_0_zero gpio1_0_one gpio1_1_tie_hi_esd gpio1_1_dm[2] gpio1_1_dm[1] gpio1_1_dm[0]
+ gpio1_1_slow gpio1_1_oe_n gpio1_1_tie_lo_esd gpio1_1_inp_dis gpio1_1_enable_vddio
+ gpio1_1_vtrip_sel gpio1_1_ib_mode_sel[1] gpio1_1_ib_mode_sel[0] gpio1_1_out gpio1_1_slew_ctl[1]
+ gpio1_1_slew_ctl[0] gpio1_1_analog_pol gpio1_1_analog_sel gpio1_1_hys_trim gpio1_0_vinref
+ gpio1_1_hld_ovr gpio1_1_in_h gpio1_1_enable_h gpio1_1_in gpio1_1_hld_h_n gpio1_1_enable_vdda_h
+ gpio1_1_analog_en gpio1_1_enable_inp_h gpio1_1_enable_vswitch_h gpio1_1_pad_a_noesd_h
+ gpio1_1_pad_a_esd_0_h gpio1_1_pad_a_esd_1_h gpio1_1_zero gpio1_1_one gpio1_2_tie_hi_esd
+ gpio1_2_dm[2] gpio1_2_dm[1] gpio1_2_dm[0] gpio1_2_slow gpio1_2_oe_n gpio1_2_tie_lo_esd
+ gpio1_2_inp_dis gpio1_2_enable_vddio gpio1_2_vtrip_sel gpio1_2_ib_mode_sel[1] gpio1_2_ib_mode_sel[0]
+ gpio1_2_out gpio1_2_slew_ctl[1] gpio1_2_slew_ctl[0] gpio1_2_analog_pol gpio1_2_analog_sel
+ gpio1_2_hys_trim gpio1_2_hld_ovr gpio1_2_in_h gpio1_2_enable_h gpio1_2_in gpio1_2_hld_h_n
+ gpio1_2_enable_vdda_h gpio1_2_analog_en gpio1_2_enable_inp_h gpio1_2_enable_vswitch_h
+ gpio1_2_pad_a_noesd_h gpio1_2_pad_a_esd_0_h gpio1_2_pad_a_esd_1_h gpio1_2_zero gpio1_2_one
+ gpio1_3_tie_hi_esd gpio1_3_dm[2] gpio1_3_dm[1] gpio1_3_dm[0] gpio1_3_slow gpio1_3_oe_n
+ gpio1_3_tie_lo_esd gpio1_3_inp_dis gpio1_3_enable_vddio gpio1_3_vtrip_sel gpio1_3_ib_mode_sel[1]
+ gpio1_3_ib_mode_sel[0] gpio1_3_out gpio1_3_slew_ctl[1] gpio1_3_slew_ctl[0] gpio1_3_analog_pol
+ gpio1_3_analog_sel gpio1_3_hys_trim gpio1_3_hld_ovr gpio1_3_in_h gpio1_3_enable_h
+ gpio1_3_in gpio1_3_hld_h_n gpio1_3_enable_vdda_h gpio1_3_analog_en gpio1_3_enable_inp_h
+ gpio1_3_enable_vswitch_h gpio1_3_pad_a_noesd_h gpio1_3_pad_a_esd_0_h gpio1_3_pad_a_esd_1_h
+ gpio1_3_zero gpio1_3_one vref_e_ref_sel[1] vref_e_ref_sel[0] vref_e_ref_sel[2] vref_e_enable_h
+ vref_e_hld_h_n vref_e_vrefgen_en vref_e_ref_sel[4] vref_e_ref_sel[3] gpio1_4_tie_hi_esd
+ gpio1_4_dm[2] gpio1_4_dm[1] gpio1_4_dm[0] gpio1_4_slow gpio1_4_oe_n gpio1_4_tie_lo_esd
+ gpio1_4_inp_dis gpio1_4_enable_vddio gpio1_4_vtrip_sel gpio1_4_ib_mode_sel[1] gpio1_4_ib_mode_sel[0]
+ gpio1_4_out gpio1_4_slew_ctl[1] gpio1_4_slew_ctl[0] gpio1_4_analog_pol gpio1_4_analog_sel
+ gpio1_4_hys_trim gpio1_4_hld_ovr gpio1_4_in_h gpio1_4_enable_h gpio1_4_in gpio1_4_hld_h_n
+ gpio1_4_enable_vdda_h gpio1_4_analog_en gpio1_4_enable_inp_h gpio1_4_enable_vswitch_h
+ gpio1_4_pad_a_noesd_h gpio1_4_pad_a_esd_0_h gpio1_4_pad_a_esd_1_h gpio1_4_zero gpio1_4_one
+ gpio1_5_tie_hi_esd gpio1_5_dm[2] gpio1_5_dm[1] gpio1_5_dm[0] gpio1_5_slow gpio1_5_oe_n
+ gpio1_5_tie_lo_esd gpio1_5_inp_dis gpio1_5_enable_vddio gpio1_5_vtrip_sel gpio1_5_ib_mode_sel[1]
+ gpio1_5_ib_mode_sel[0] gpio1_5_out gpio1_5_slew_ctl[1] gpio1_5_slew_ctl[0] gpio1_5_analog_pol
+ gpio1_5_analog_sel gpio1_5_hys_trim gpio1_5_hld_ovr gpio1_5_in_h gpio1_5_enable_h
+ gpio1_5_in gpio1_5_hld_h_n gpio1_5_enable_vdda_h gpio1_5_analog_en gpio1_5_enable_inp_h
+ gpio1_5_enable_vswitch_h gpio1_5_pad_a_noesd_h gpio1_5_pad_a_esd_0_h gpio1_5_pad_a_esd_1_h
+ gpio1_5_zero gpio1_5_one gpio1_6_tie_hi_esd gpio1_6_dm[2] gpio1_6_dm[1] gpio1_6_dm[0]
+ gpio1_6_slow gpio1_6_oe_n gpio1_6_tie_lo_esd gpio1_6_inp_dis gpio1_6_enable_vddio
+ gpio1_6_vtrip_sel gpio1_6_ib_mode_sel[1] gpio1_6_ib_mode_sel[0] gpio1_6_out gpio1_6_slew_ctl[1]
+ gpio1_6_slew_ctl[0] gpio1_6_analog_pol gpio1_6_analog_sel gpio1_6_hys_trim gpio1_6_hld_ovr
+ gpio1_6_in_h gpio1_6_enable_h gpio1_6_in gpio1_6_hld_h_n gpio1_6_enable_vdda_h gpio1_6_analog_en
+ gpio1_6_enable_inp_h gpio1_6_enable_vswitch_h gpio1_6_pad_a_noesd_h gpio1_6_pad_a_esd_0_h
+ gpio1_6_pad_a_esd_1_h gpio1_6_zero gpio1_6_one gpio1_7_tie_hi_esd gpio1_7_dm[2]
+ gpio1_7_dm[1] gpio1_7_dm[0] gpio1_7_slow gpio1_7_oe_n gpio1_7_tie_lo_esd gpio1_7_inp_dis
+ gpio1_7_enable_vddio gpio1_7_vtrip_sel gpio1_7_ib_mode_sel[1] gpio1_7_ib_mode_sel[0]
+ gpio1_7_out gpio1_7_slew_ctl[1] gpio1_7_slew_ctl[0] gpio1_7_analog_pol gpio1_7_analog_sel
+ gpio1_7_hys_trim vcap_e_cpos gpio1_7_hld_ovr gpio1_7_in_h gpio1_7_enable_h gpio1_7_in
+ gpio1_7_hld_h_n gpio1_7_enable_vdda_h gpio1_7_analog_en gpio1_7_enable_inp_h gpio1_7_enable_vswitch_h
+ gpio1_7_pad_a_noesd_h gpio1_7_pad_a_esd_0_h gpio1_7_pad_a_esd_1_h gpio1_7_zero gpio1_7_one
+ gpio2_0_tie_lo_esd gpio2_0_in gpio2_0_tie_hi_esd gpio2_0_enable_vddio gpio2_0_slow
+ gpio2_0_pad_a_esd_0_h gpio2_0_pad_a_esd_1_h gpio2_0_pad_a_noesd_h gpio2_0_analog_en
+ gpio2_0_analog_pol gpio2_0_inp_dis gpio2_0_enable_inp_h gpio2_0_enable_h gpio2_0_hld_h_n
+ gpio2_0_analog_sel gpio2_0_dm[2] gpio2_0_dm[1] gpio2_0_dm[0] gpio2_0_hld_ovr gpio2_0_out
+ gpio2_0_enable_vswitch_h gpio2_0_enable_vdda_h gpio2_0_vtrip_sel gpio2_0_ib_mode_sel
+ gpio2_0_oe_n gpio2_0_in_h gpio2_0_zero gpio2_0_one gpio2_1_tie_lo_esd gpio2_1_in
+ gpio2_1_tie_hi_esd gpio2_1_enable_vddio gpio2_1_slow gpio2_1_pad_a_esd_0_h gpio2_1_pad_a_esd_1_h
+ gpio2_1_pad_a_noesd_h gpio2_1_analog_en gpio2_1_analog_pol gpio2_1_inp_dis gpio2_1_enable_inp_h
+ gpio2_1_enable_h gpio2_1_hld_h_n gpio2_1_analog_sel gpio2_1_dm[2] gpio2_1_dm[1]
+ gpio2_1_dm[0] gpio2_1_hld_ovr gpio2_1_out gpio2_1_enable_vswitch_h gpio2_1_enable_vdda_h
+ gpio2_1_vtrip_sel gpio2_1_ib_mode_sel gpio2_1_oe_n gpio2_1_in_h gpio2_1_zero gpio2_1_one
+ gpio2_2_tie_lo_esd gpio2_2_in gpio2_2_tie_hi_esd gpio2_2_enable_vddio gpio2_2_slow
+ gpio2_2_pad_a_esd_0_h gpio2_2_pad_a_esd_1_h gpio2_2_pad_a_noesd_h gpio2_2_analog_en
+ gpio2_2_analog_pol gpio2_2_inp_dis gpio2_2_enable_inp_h gpio2_2_enable_h gpio2_2_hld_h_n
+ gpio2_2_analog_sel gpio2_2_dm[2] gpio2_2_dm[1] gpio2_2_dm[0] gpio2_2_hld_ovr gpio2_2_out
+ gpio2_2_enable_vswitch_h gpio2_2_enable_vdda_h gpio2_2_vtrip_sel gpio2_2_ib_mode_sel
+ gpio2_2_oe_n gpio2_2_in_h gpio2_2_zero gpio2_2_one gpio2_3_tie_lo_esd gpio2_3_in
+ gpio2_3_tie_hi_esd gpio2_3_enable_vddio gpio2_3_slow gpio2_3_pad_a_esd_0_h gpio2_3_pad_a_esd_1_h
+ gpio2_3_pad_a_noesd_h gpio2_3_analog_en gpio2_3_analog_pol gpio2_3_inp_dis gpio2_3_enable_inp_h
+ gpio2_3_enable_h gpio2_3_hld_h_n gpio2_3_analog_sel gpio2_3_dm[2] gpio2_3_dm[1]
+ gpio2_3_dm[0] gpio2_3_hld_ovr gpio2_3_out gpio2_3_enable_vswitch_h gpio2_3_enable_vdda_h
+ gpio2_3_vtrip_sel gpio2_3_ib_mode_sel gpio2_3_oe_n gpio2_3_in_h gpio2_3_zero gpio2_3_one
+ gpio2_4_tie_lo_esd gpio2_4_in gpio2_4_tie_hi_esd gpio2_4_enable_vddio gpio2_4_slow
+ gpio2_4_pad_a_esd_0_h gpio2_4_pad_a_esd_1_h gpio2_4_pad_a_noesd_h gpio2_4_analog_en
+ gpio2_4_analog_pol gpio2_4_inp_dis gpio2_4_enable_inp_h gpio2_4_enable_h gpio2_4_hld_h_n
+ gpio2_4_analog_sel gpio2_4_dm[2] gpio2_4_dm[1] gpio2_4_dm[0] gpio2_4_hld_ovr gpio2_4_out
+ gpio2_4_enable_vswitch_h gpio2_4_enable_vdda_h gpio2_4_vtrip_sel gpio2_4_ib_mode_sel
+ gpio2_4_oe_n gpio2_4_in_h gpio2_4_zero gpio2_4_one gpio2_5_tie_lo_esd gpio2_5_in
+ gpio2_5_tie_hi_esd gpio2_5_enable_vddio gpio2_5_slow gpio2_5_pad_a_esd_0_h gpio2_5_pad_a_esd_1_h
+ gpio2_5_pad_a_noesd_h gpio2_5_analog_en gpio2_5_analog_pol gpio2_5_inp_dis gpio2_5_enable_inp_h
+ gpio2_5_enable_h gpio2_5_hld_h_n gpio2_5_analog_sel gpio2_5_dm[2] gpio2_5_dm[1]
+ gpio2_5_dm[0] gpio2_5_hld_ovr gpio2_5_out gpio2_5_enable_vswitch_h gpio2_5_enable_vdda_h
+ gpio2_5_vtrip_sel gpio2_5_ib_mode_sel gpio2_5_oe_n gpio2_5_in_h gpio2_5_zero gpio2_5_one
+ gpio2_6_tie_lo_esd gpio2_6_in gpio2_6_tie_hi_esd gpio2_6_enable_vddio gpio2_6_slow
+ gpio2_6_pad_a_esd_0_h gpio2_6_pad_a_esd_1_h gpio2_6_pad_a_noesd_h gpio2_6_analog_en
+ gpio2_6_analog_pol gpio2_6_inp_dis gpio2_6_enable_inp_h gpio2_6_enable_h gpio2_6_hld_h_n
+ gpio2_6_analog_sel gpio2_6_dm[2] gpio2_6_dm[1] gpio2_6_dm[0] gpio2_6_hld_ovr gpio2_6_out
+ gpio2_6_enable_vswitch_h gpio2_6_enable_vdda_h gpio2_6_vtrip_sel gpio2_6_ib_mode_sel
+ gpio2_6_oe_n gpio2_6_in_h gpio2_6_zero gpio2_6_one gpio2_7_tie_lo_esd gpio2_7_in
+ gpio2_7_tie_hi_esd gpio2_7_enable_vddio gpio2_7_slow gpio2_7_pad_a_esd_0_h gpio2_7_pad_a_esd_1_h
+ gpio2_7_pad_a_noesd_h gpio2_7_analog_en gpio2_7_analog_pol gpio2_7_inp_dis gpio2_7_enable_inp_h
+ gpio2_7_enable_h gpio2_7_hld_h_n gpio2_7_analog_sel gpio2_7_dm[2] gpio2_7_dm[1]
+ gpio2_7_dm[0] gpio2_7_hld_ovr gpio2_7_out gpio2_7_enable_vswitch_h gpio2_7_enable_vdda_h
+ gpio2_7_vtrip_sel gpio2_7_ib_mode_sel gpio2_7_oe_n gpio2_7_in_h gpio2_7_zero gpio2_7_one
+ muxsplit_ne_hld_vdda_h_n muxsplit_ne_enable_vdda_h muxsplit_ne_switch_aa_sl muxsplit_ne_switch_aa_s0
+ muxsplit_ne_switch_bb_s0 muxsplit_ne_switch_bb_sl muxsplit_ne_switch_bb_sr muxsplit_ne_switch_aa_sr
+ gpio3_0_tie_lo_esd gpio3_0_in gpio3_0_tie_hi_esd gpio3_0_enable_vddio gpio3_0_slow
+ gpio3_0_pad_a_esd_0_h gpio3_0_pad_a_esd_1_h gpio3_0_pad_a_noesd_h gpio3_0_analog_en
+ gpio3_0_analog_pol gpio3_0_inp_dis gpio3_0_enable_inp_h gpio3_0_enable_h gpio3_0_hld_h_n
+ gpio3_0_analog_sel gpio3_0_dm[2] gpio3_0_dm[1] gpio3_0_dm[0] gpio3_0_hld_ovr gpio3_0_out
+ gpio3_0_enable_vswitch_h gpio3_0_enable_vdda_h gpio3_0_vtrip_sel gpio3_0_ib_mode_sel
+ gpio3_0_oe_n gpio3_0_in_h gpio3_0_zero gpio3_0_one gpio3_1_tie_lo_esd gpio3_1_in
+ gpio3_1_tie_hi_esd gpio3_1_enable_vddio gpio3_1_slow gpio3_1_pad_a_esd_0_h gpio3_1_pad_a_esd_1_h
+ gpio3_1_pad_a_noesd_h gpio3_1_analog_en gpio3_1_analog_pol gpio3_1_inp_dis gpio3_1_enable_inp_h
+ gpio3_1_enable_h gpio3_1_hld_h_n gpio3_1_analog_sel gpio3_1_dm[2] gpio3_1_dm[1]
+ gpio3_1_dm[0] gpio3_1_hld_ovr gpio3_1_out gpio3_1_enable_vswitch_h gpio3_1_enable_vdda_h
+ gpio3_1_vtrip_sel gpio3_1_ib_mode_sel gpio3_1_oe_n gpio3_1_in_h gpio3_1_zero gpio3_1_one
+ gpio3_2_tie_lo_esd gpio3_2_in gpio3_2_tie_hi_esd gpio3_2_enable_vddio gpio3_2_slow
+ gpio3_2_pad_a_esd_0_h gpio3_2_pad_a_esd_1_h gpio3_2_pad_a_noesd_h gpio3_2_analog_en
+ gpio3_2_analog_pol gpio3_2_inp_dis gpio3_2_enable_inp_h gpio3_2_enable_h gpio3_2_hld_h_n
+ gpio3_2_analog_sel gpio3_2_dm[2] gpio3_2_dm[1] gpio3_2_dm[0] gpio3_2_hld_ovr gpio3_2_out
+ gpio3_2_enable_vswitch_h gpio3_2_enable_vdda_h gpio3_2_vtrip_sel gpio3_2_ib_mode_sel
+ gpio3_2_oe_n gpio3_2_in_h gpio3_2_zero gpio3_2_one gpio3_3_tie_lo_esd gpio3_3_in
+ gpio3_3_tie_hi_esd gpio3_3_enable_vddio gpio3_3_slow gpio3_3_pad_a_esd_0_h gpio3_3_pad_a_esd_1_h
+ gpio3_3_pad_a_noesd_h gpio3_3_analog_en gpio3_3_analog_pol gpio3_3_inp_dis gpio3_3_enable_inp_h
+ gpio3_3_enable_h gpio3_3_hld_h_n gpio3_3_analog_sel gpio3_3_dm[2] gpio3_3_dm[1]
+ gpio3_3_dm[0] gpio3_3_hld_ovr gpio3_3_out gpio3_3_enable_vswitch_h gpio3_3_enable_vdda_h
+ gpio3_3_vtrip_sel gpio3_3_ib_mode_sel gpio3_3_oe_n gpio3_3_in_h gpio3_3_zero gpio3_3_one
+ gpio3_4_tie_lo_esd gpio3_4_in gpio3_4_tie_hi_esd gpio3_4_enable_vddio gpio3_4_slow
+ gpio3_4_pad_a_esd_0_h gpio3_4_pad_a_esd_1_h gpio3_4_pad_a_noesd_h gpio3_4_analog_en
+ gpio3_4_analog_pol gpio3_4_inp_dis gpio3_4_enable_inp_h gpio3_4_enable_h gpio3_4_hld_h_n
+ gpio3_4_analog_sel gpio3_4_dm[2] gpio3_4_dm[1] gpio3_4_dm[0] gpio3_4_hld_ovr gpio3_4_out
+ gpio3_4_enable_vswitch_h gpio3_4_enable_vdda_h gpio3_4_vtrip_sel gpio3_4_ib_mode_sel
+ gpio3_4_oe_n gpio3_4_in_h gpio3_4_zero gpio3_4_one gpio3_5_tie_lo_esd gpio3_5_in
+ gpio3_5_tie_hi_esd gpio3_5_enable_vddio gpio3_5_slow gpio3_5_pad_a_esd_0_h gpio3_5_pad_a_esd_1_h
+ gpio3_5_pad_a_noesd_h gpio3_5_analog_en gpio3_5_analog_pol gpio3_5_inp_dis gpio3_5_enable_inp_h
+ gpio3_5_enable_h gpio3_5_hld_h_n gpio3_5_analog_sel gpio3_5_dm[2] gpio3_5_dm[1]
+ gpio3_5_dm[0] gpio3_5_hld_ovr gpio3_5_out gpio3_5_enable_vswitch_h gpio3_5_enable_vdda_h
+ gpio3_5_vtrip_sel gpio3_5_ib_mode_sel gpio3_5_oe_n gpio3_5_in_h gpio3_5_zero gpio3_5_one
+ gpio3_6_tie_lo_esd gpio3_6_in gpio3_6_tie_hi_esd gpio3_6_enable_vddio gpio3_6_slow
+ gpio3_6_pad_a_esd_0_h gpio3_6_pad_a_esd_1_h gpio3_6_pad_a_noesd_h gpio3_6_analog_en
+ gpio3_6_analog_pol gpio3_6_inp_dis gpio3_6_enable_inp_h gpio3_6_enable_h gpio3_6_hld_h_n
+ gpio3_6_analog_sel gpio3_6_dm[2] gpio3_6_dm[1] gpio3_6_dm[0] gpio3_6_hld_ovr gpio3_6_out
+ gpio3_6_enable_vswitch_h gpio3_6_enable_vdda_h gpio3_6_vtrip_sel gpio3_6_ib_mode_sel
+ gpio3_6_oe_n gpio3_6_in_h gpio3_6_zero gpio3_6_one gpio3_7_tie_lo_esd gpio3_7_in
+ gpio3_7_tie_hi_esd gpio3_7_enable_vddio gpio3_7_slow gpio3_7_pad_a_esd_0_h gpio3_7_pad_a_esd_1_h
+ gpio3_7_pad_a_noesd_h gpio3_7_analog_en gpio3_7_analog_pol gpio3_7_inp_dis gpio3_7_enable_inp_h
+ gpio3_7_enable_h gpio3_7_hld_h_n gpio3_7_analog_sel gpio3_7_dm[2] gpio3_7_dm[1]
+ gpio3_7_dm[0] gpio3_7_hld_ovr gpio3_7_out gpio3_7_enable_vswitch_h gpio3_7_enable_vdda_h
+ gpio3_7_vtrip_sel gpio3_7_ib_mode_sel gpio3_7_oe_n gpio3_7_in_h gpio3_7_zero gpio3_7_one
+ analog_0_core analog_1_core gpio4_0_tie_lo_esd gpio4_0_in gpio4_0_tie_hi_esd gpio4_0_enable_vddio
+ gpio4_0_slow gpio4_0_pad_a_esd_0_h gpio4_0_pad_a_esd_1_h gpio4_0_pad_a_noesd_h gpio4_0_analog_en
+ gpio4_0_analog_pol gpio4_0_inp_dis gpio4_0_enable_inp_h gpio4_0_enable_h gpio4_0_hld_h_n
+ gpio4_0_analog_sel gpio4_0_dm[2] gpio4_0_dm[1] gpio4_0_dm[0] gpio4_0_hld_ovr gpio4_0_out
+ gpio4_0_enable_vswitch_h gpio4_0_enable_vdda_h gpio4_0_vtrip_sel gpio4_0_ib_mode_sel
+ gpio4_0_oe_n gpio4_0_in_h gpio4_0_zero gpio4_0_one gpio4_1_tie_lo_esd gpio4_1_in
+ gpio4_1_tie_hi_esd gpio4_1_enable_vddio gpio4_1_slow gpio4_1_pad_a_esd_0_h gpio4_1_pad_a_esd_1_h
+ gpio4_1_pad_a_noesd_h gpio4_1_analog_en gpio4_1_analog_pol gpio4_1_inp_dis gpio4_1_enable_inp_h
+ gpio4_1_enable_h gpio4_1_hld_h_n gpio4_1_analog_sel gpio4_1_dm[2] gpio4_1_dm[1]
+ gpio4_1_dm[0] gpio4_1_hld_ovr gpio4_1_out gpio4_1_enable_vswitch_h gpio4_1_enable_vdda_h
+ gpio4_1_vtrip_sel gpio4_1_ib_mode_sel gpio4_1_oe_n gpio4_1_in_h gpio4_1_zero gpio4_1_one
+ gpio4_2_tie_lo_esd gpio4_2_in gpio4_2_tie_hi_esd gpio4_2_enable_vddio gpio4_2_slow
+ gpio4_2_pad_a_esd_0_h gpio4_2_pad_a_esd_1_h gpio4_2_pad_a_noesd_h gpio4_2_analog_en
+ gpio4_2_analog_pol gpio4_2_inp_dis gpio4_2_enable_inp_h gpio4_2_enable_h gpio4_2_hld_h_n
+ gpio4_2_analog_sel gpio4_2_dm[2] gpio4_2_dm[1] gpio4_2_dm[0] gpio4_2_hld_ovr gpio4_2_out
+ gpio4_2_enable_vswitch_h gpio4_2_enable_vdda_h gpio4_2_vtrip_sel gpio4_2_ib_mode_sel
+ gpio4_2_oe_n gpio4_2_in_h gpio4_2_zero gpio4_2_one gpio4_3_tie_lo_esd gpio4_3_in
+ gpio4_3_tie_hi_esd gpio4_3_enable_vddio gpio4_3_slow gpio4_3_pad_a_esd_0_h gpio4_3_pad_a_esd_1_h
+ gpio4_3_pad_a_noesd_h gpio4_3_analog_en gpio4_3_analog_pol gpio4_3_inp_dis gpio4_3_enable_inp_h
+ gpio4_3_enable_h gpio4_3_hld_h_n gpio4_3_analog_sel gpio4_3_dm[2] gpio4_3_dm[1]
+ gpio4_3_dm[0] gpio4_3_hld_ovr gpio4_3_out gpio4_3_enable_vswitch_h gpio4_3_enable_vdda_h
+ gpio4_3_vtrip_sel gpio4_3_ib_mode_sel gpio4_3_oe_n gpio4_3_in_h gpio4_3_zero gpio4_3_one
+ gpio4_4_tie_lo_esd gpio4_4_in gpio4_4_tie_hi_esd gpio4_4_enable_vddio gpio4_4_slow
+ gpio4_4_pad_a_esd_0_h gpio4_4_pad_a_esd_1_h gpio4_4_pad_a_noesd_h gpio4_4_analog_en
+ gpio4_4_analog_pol gpio4_4_inp_dis gpio4_4_enable_inp_h gpio4_4_enable_h gpio4_4_hld_h_n
+ gpio4_4_analog_sel gpio4_4_dm[2] gpio4_4_dm[1] gpio4_4_dm[0] gpio4_4_hld_ovr gpio4_4_out
+ gpio4_4_enable_vswitch_h gpio4_4_enable_vdda_h gpio4_4_vtrip_sel gpio4_4_ib_mode_sel
+ gpio4_4_oe_n gpio4_4_in_h gpio4_4_zero gpio4_4_one gpio4_5_tie_lo_esd gpio4_5_in
+ gpio4_5_tie_hi_esd gpio4_5_enable_vddio gpio4_5_slow gpio4_5_pad_a_esd_0_h gpio4_5_pad_a_esd_1_h
+ gpio4_5_pad_a_noesd_h gpio4_5_analog_en gpio4_5_analog_pol gpio4_5_inp_dis gpio4_5_enable_inp_h
+ gpio4_5_enable_h gpio4_5_hld_h_n gpio4_5_analog_sel gpio4_5_dm[2] gpio4_5_dm[1]
+ gpio4_5_dm[0] gpio4_5_hld_ovr gpio4_5_out gpio4_5_enable_vswitch_h gpio4_5_enable_vdda_h
+ gpio4_5_vtrip_sel gpio4_5_ib_mode_sel gpio4_5_oe_n gpio4_5_in_h gpio4_5_zero gpio4_5_one
+ gpio4_6_tie_lo_esd gpio4_6_in gpio4_6_tie_hi_esd gpio4_6_enable_vddio gpio4_6_slow
+ gpio4_6_pad_a_esd_0_h gpio4_6_pad_a_esd_1_h gpio4_6_pad_a_noesd_h gpio4_6_analog_en
+ gpio4_6_analog_pol gpio4_6_inp_dis gpio4_6_enable_inp_h gpio4_6_enable_h gpio4_6_hld_h_n
+ gpio4_6_analog_sel gpio4_6_dm[2] gpio4_6_dm[1] gpio4_6_dm[0] gpio4_6_hld_ovr gpio4_6_out
+ gpio4_6_enable_vswitch_h gpio4_6_enable_vdda_h gpio4_6_vtrip_sel gpio4_6_ib_mode_sel
+ gpio4_6_oe_n gpio4_6_in_h gpio4_6_zero gpio4_6_one gpio4_7_tie_lo_esd gpio4_7_in
+ gpio4_7_tie_hi_esd gpio4_7_enable_vddio gpio4_7_slow gpio4_7_pad_a_esd_0_h gpio4_7_pad_a_esd_1_h
+ gpio4_7_pad_a_noesd_h gpio4_7_analog_en gpio4_7_analog_pol gpio4_7_inp_dis gpio4_7_enable_inp_h
+ gpio4_7_enable_h gpio4_7_hld_h_n gpio4_7_analog_sel gpio4_7_dm[2] gpio4_7_dm[1]
+ gpio4_7_dm[0] gpio4_7_hld_ovr gpio4_7_out gpio4_7_enable_vswitch_h gpio4_7_enable_vdda_h
+ gpio4_7_vtrip_sel gpio4_7_ib_mode_sel gpio4_7_oe_n gpio4_7_in_h gpio4_7_zero gpio4_7_one
+ muxsplit_nw_hld_vdda_h_n muxsplit_nw_enable_vdda_h muxsplit_nw_switch_aa_sl muxsplit_nw_switch_aa_s0
+ muxsplit_nw_switch_bb_s0 muxsplit_nw_switch_bb_sl muxsplit_nw_switch_bb_sr muxsplit_nw_switch_aa_sr
+ gpio5_0_tie_lo_esd gpio5_0_in gpio5_0_tie_hi_esd gpio5_0_enable_vddio gpio5_0_slow
+ gpio5_0_pad_a_esd_0_h gpio5_0_pad_a_esd_1_h gpio5_0_pad_a_noesd_h gpio5_0_analog_en
+ gpio5_0_analog_pol gpio5_0_inp_dis gpio5_0_enable_inp_h gpio5_0_enable_h gpio5_0_hld_h_n
+ gpio5_0_analog_sel gpio5_0_dm[2] gpio5_0_dm[1] gpio5_0_dm[0] gpio5_0_hld_ovr gpio5_0_out
+ gpio5_0_enable_vswitch_h gpio5_0_enable_vdda_h gpio5_0_vtrip_sel gpio5_0_ib_mode_sel
+ gpio5_0_oe_n gpio5_0_in_h gpio5_0_zero gpio5_0_one gpio5_1_tie_lo_esd gpio5_1_in
+ gpio5_1_tie_hi_esd gpio5_1_enable_vddio gpio5_1_slow gpio5_1_pad_a_esd_0_h gpio5_1_pad_a_esd_1_h
+ gpio5_1_pad_a_noesd_h gpio5_1_analog_en gpio5_1_analog_pol gpio5_1_inp_dis gpio5_1_enable_inp_h
+ gpio5_1_enable_h gpio5_1_hld_h_n gpio5_1_analog_sel gpio5_1_dm[2] gpio5_1_dm[1]
+ gpio5_1_dm[0] gpio5_1_hld_ovr gpio5_1_out gpio5_1_enable_vswitch_h gpio5_1_enable_vdda_h
+ gpio5_1_vtrip_sel gpio5_1_ib_mode_sel gpio5_1_oe_n gpio5_1_in_h gpio5_1_zero gpio5_1_one
+ gpio5_2_tie_lo_esd gpio5_2_in gpio5_2_tie_hi_esd gpio5_2_enable_vddio gpio5_2_slow
+ gpio5_2_pad_a_esd_0_h gpio5_2_pad_a_esd_1_h gpio5_2_pad_a_noesd_h gpio5_2_analog_en
+ gpio5_2_analog_pol gpio5_2_inp_dis gpio5_2_enable_inp_h gpio5_2_enable_h gpio5_2_hld_h_n
+ gpio5_2_analog_sel gpio5_2_dm[2] gpio5_2_dm[1] gpio5_2_dm[0] gpio5_2_hld_ovr gpio5_2_out
+ gpio5_2_enable_vswitch_h gpio5_2_enable_vdda_h gpio5_2_vtrip_sel gpio5_2_ib_mode_sel
+ gpio5_2_oe_n gpio5_2_in_h gpio5_2_zero gpio5_2_one gpio5_3_tie_lo_esd gpio5_3_in
+ gpio5_3_tie_hi_esd gpio5_3_enable_vddio gpio5_3_slow gpio5_3_pad_a_esd_0_h gpio5_3_pad_a_esd_1_h
+ gpio5_3_pad_a_noesd_h gpio5_3_analog_en gpio5_3_analog_pol gpio5_3_inp_dis gpio5_3_enable_inp_h
+ gpio5_3_enable_h gpio5_3_hld_h_n gpio5_3_analog_sel gpio5_3_dm[2] gpio5_3_dm[1]
+ gpio5_3_dm[0] gpio5_3_hld_ovr gpio5_3_out gpio5_3_enable_vswitch_h gpio5_3_enable_vdda_h
+ gpio5_3_vtrip_sel gpio5_3_ib_mode_sel gpio5_3_oe_n gpio5_3_in_h gpio5_3_zero gpio5_3_one
+ gpio5_4_tie_lo_esd gpio5_4_in gpio5_4_tie_hi_esd gpio5_4_enable_vddio gpio5_4_slow
+ gpio5_4_pad_a_esd_0_h gpio5_4_pad_a_esd_1_h gpio5_4_pad_a_noesd_h gpio5_4_analog_en
+ gpio5_4_analog_pol gpio5_4_inp_dis gpio5_4_enable_inp_h gpio5_4_enable_h gpio5_4_hld_h_n
+ gpio5_4_analog_sel gpio5_4_dm[2] gpio5_4_dm[1] gpio5_4_dm[0] gpio5_4_hld_ovr gpio5_4_out
+ gpio5_4_enable_vswitch_h gpio5_4_enable_vdda_h gpio5_4_vtrip_sel gpio5_4_ib_mode_sel
+ gpio5_4_oe_n gpio5_4_in_h gpio5_4_zero gpio5_4_one gpio5_5_tie_lo_esd gpio5_5_in
+ gpio5_5_tie_hi_esd gpio5_5_enable_vddio gpio5_5_slow gpio5_5_pad_a_esd_0_h gpio5_5_pad_a_esd_1_h
+ gpio5_5_pad_a_noesd_h gpio5_5_analog_en gpio5_5_analog_pol gpio5_5_inp_dis gpio5_5_enable_inp_h
+ gpio5_5_enable_h gpio5_5_hld_h_n gpio5_5_analog_sel gpio5_5_dm[2] gpio5_5_dm[1]
+ gpio5_5_dm[0] gpio5_5_hld_ovr gpio5_5_out gpio5_5_enable_vswitch_h gpio5_5_enable_vdda_h
+ gpio5_5_vtrip_sel gpio5_5_ib_mode_sel gpio5_5_oe_n gpio5_5_in_h gpio5_5_zero gpio5_5_one
+ gpio5_6_tie_lo_esd gpio5_6_in gpio5_6_tie_hi_esd gpio5_6_enable_vddio gpio5_6_slow
+ gpio5_6_pad_a_esd_0_h gpio5_6_pad_a_esd_1_h gpio5_6_pad_a_noesd_h gpio5_6_analog_en
+ gpio5_6_analog_pol gpio5_6_inp_dis gpio5_6_enable_inp_h gpio5_6_enable_h gpio5_6_hld_h_n
+ gpio5_6_analog_sel gpio5_6_dm[2] gpio5_6_dm[1] gpio5_6_dm[0] gpio5_6_hld_ovr gpio5_6_out
+ gpio5_6_enable_vswitch_h gpio5_6_enable_vdda_h gpio5_6_vtrip_sel gpio5_6_ib_mode_sel
+ gpio5_6_oe_n gpio5_6_in_h gpio5_6_zero gpio5_6_one gpio5_7_tie_lo_esd gpio5_7_in
+ gpio5_7_tie_hi_esd gpio5_7_enable_vddio gpio5_7_slow gpio5_7_pad_a_esd_0_h gpio5_7_pad_a_esd_1_h
+ gpio5_7_pad_a_noesd_h gpio5_7_analog_en gpio5_7_analog_pol gpio5_7_inp_dis gpio5_7_enable_inp_h
+ gpio5_7_enable_h gpio5_7_hld_h_n gpio5_7_analog_sel gpio5_7_dm[2] gpio5_7_dm[1]
+ gpio5_7_dm[0] gpio5_7_hld_ovr gpio5_7_out gpio5_7_enable_vswitch_h gpio5_7_enable_vdda_h
+ gpio5_7_vtrip_sel gpio5_7_ib_mode_sel gpio5_7_oe_n gpio5_7_in_h gpio5_7_zero gpio5_7_one
+ gpio6_0_tie_hi_esd gpio6_0_dm[2] gpio6_0_dm[1] gpio6_0_dm[0] gpio6_0_slow gpio6_0_oe_n
+ gpio6_0_tie_lo_esd gpio6_0_inp_dis gpio6_0_enable_vddio gpio6_0_vtrip_sel gpio6_0_ib_mode_sel[1]
+ gpio6_0_ib_mode_sel[0] gpio6_0_out gpio6_0_slew_ctl[1] gpio6_0_slew_ctl[0] gpio6_0_analog_pol
+ gpio6_0_analog_sel gpio6_0_hys_trim vcap_w_cpos gpio6_0_hld_ovr gpio6_0_in_h gpio6_0_enable_h
+ gpio6_0_in gpio6_0_hld_h_n gpio6_0_enable_vdda_h gpio6_0_analog_en gpio6_0_enable_inp_h
+ gpio6_0_enable_vswitch_h gpio6_0_pad_a_noesd_h gpio6_0_pad_a_esd_0_h gpio6_0_pad_a_esd_1_h
+ gpio6_0_zero gpio6_0_one gpio6_1_tie_hi_esd gpio6_1_dm[2] gpio6_1_dm[1] gpio6_1_dm[0]
+ gpio6_1_slow gpio6_1_oe_n gpio6_1_tie_lo_esd gpio6_1_inp_dis gpio6_1_enable_vddio
+ gpio6_1_vtrip_sel gpio6_1_ib_mode_sel[1] gpio6_1_ib_mode_sel[0] gpio6_1_out gpio6_1_slew_ctl[1]
+ gpio6_1_slew_ctl[0] gpio6_1_analog_pol gpio6_1_analog_sel gpio6_1_hys_trim gpio6_1_hld_ovr
+ gpio6_1_in_h gpio6_1_enable_h gpio6_1_in gpio6_1_hld_h_n gpio6_1_enable_vdda_h gpio6_1_analog_en
+ gpio6_1_enable_inp_h gpio6_1_enable_vswitch_h gpio6_1_pad_a_noesd_h gpio6_1_pad_a_esd_0_h
+ gpio6_1_pad_a_esd_1_h gpio6_1_zero gpio6_1_one gpio6_2_tie_hi_esd gpio6_2_dm[2]
+ gpio6_2_dm[1] gpio6_2_dm[0] gpio6_2_slow gpio6_2_oe_n gpio6_2_tie_lo_esd gpio6_2_inp_dis
+ gpio6_2_enable_vddio gpio6_2_vtrip_sel gpio6_2_ib_mode_sel[1] gpio6_2_ib_mode_sel[0]
+ gpio6_2_out gpio6_2_slew_ctl[1] gpio6_2_slew_ctl[0] gpio6_2_analog_pol gpio6_2_analog_sel
+ gpio6_2_hys_trim gpio6_2_hld_ovr gpio6_2_in_h gpio6_2_enable_h gpio6_2_in gpio6_2_hld_h_n
+ gpio6_2_enable_vdda_h gpio6_2_analog_en gpio6_2_enable_inp_h gpio6_2_enable_vswitch_h
+ gpio6_2_pad_a_noesd_h gpio6_2_pad_a_esd_0_h gpio6_2_pad_a_esd_1_h gpio6_2_zero gpio6_2_one
+ gpio6_3_tie_hi_esd gpio6_3_dm[2] gpio6_3_dm[1] gpio6_3_dm[0] gpio6_3_slow gpio6_3_oe_n
+ gpio6_3_tie_lo_esd gpio6_3_inp_dis gpio6_3_enable_vddio gpio6_3_vtrip_sel gpio6_3_ib_mode_sel[1]
+ gpio6_3_ib_mode_sel[0] gpio6_3_out gpio6_3_slew_ctl[1] gpio6_3_slew_ctl[0] gpio6_3_analog_pol
+ gpio6_3_analog_sel gpio6_3_hys_trim gpio6_3_hld_ovr gpio6_3_in_h gpio6_3_enable_h
+ gpio6_3_in gpio6_3_hld_h_n gpio6_3_enable_vdda_h gpio6_3_analog_en gpio6_3_enable_inp_h
+ gpio6_3_enable_vswitch_h gpio6_3_pad_a_noesd_h gpio6_3_pad_a_esd_0_h gpio6_3_pad_a_esd_1_h
+ gpio6_3_zero gpio6_3_one vref_w_ref_sel[1] vref_w_ref_sel[0] vref_w_ref_sel[2] vref_w_enable_h
+ vref_w_hld_h_n vref_w_vrefgen_en vref_w_ref_sel[4] vref_w_ref_sel[3] gpio6_4_tie_hi_esd
+ gpio6_4_dm[2] gpio6_4_dm[1] gpio6_4_dm[0] gpio6_4_slow gpio6_4_oe_n gpio6_4_tie_lo_esd
+ gpio6_4_inp_dis gpio6_4_enable_vddio gpio6_4_vtrip_sel gpio6_4_ib_mode_sel[1] gpio6_4_ib_mode_sel[0]
+ gpio6_4_out gpio6_4_slew_ctl[1] gpio6_4_slew_ctl[0] gpio6_4_analog_pol gpio6_4_analog_sel
+ gpio6_4_hys_trim gpio6_7_vinref gpio6_4_hld_ovr gpio6_4_in_h gpio6_4_enable_h gpio6_4_in
+ gpio6_4_hld_h_n gpio6_4_enable_vdda_h gpio6_4_analog_en gpio6_4_enable_inp_h gpio6_4_enable_vswitch_h
+ gpio6_4_pad_a_noesd_h gpio6_4_pad_a_esd_0_h gpio6_4_pad_a_esd_1_h gpio6_4_zero gpio6_4_one
+ gpio6_5_tie_hi_esd gpio6_5_dm[2] gpio6_5_dm[1] gpio6_5_dm[0] gpio6_5_slow gpio6_5_oe_n
+ gpio6_5_tie_lo_esd gpio6_5_inp_dis gpio6_5_enable_vddio gpio6_5_vtrip_sel gpio6_5_ib_mode_sel[1]
+ gpio6_5_ib_mode_sel[0] gpio6_5_out gpio6_5_slew_ctl[1] gpio6_5_slew_ctl[0] gpio6_5_analog_pol
+ gpio6_5_analog_sel gpio6_5_hys_trim gpio6_5_hld_ovr gpio6_5_in_h gpio6_5_enable_h
+ gpio6_5_in gpio6_5_hld_h_n gpio6_5_enable_vdda_h gpio6_5_analog_en gpio6_5_enable_inp_h
+ gpio6_5_enable_vswitch_h gpio6_5_pad_a_noesd_h gpio6_5_pad_a_esd_0_h gpio6_5_pad_a_esd_1_h
+ gpio6_5_zero gpio6_5_one gpio6_6_tie_hi_esd gpio6_6_dm[2] gpio6_6_dm[1] gpio6_6_dm[0]
+ gpio6_6_slow gpio6_6_oe_n gpio6_6_tie_lo_esd gpio6_6_inp_dis gpio6_6_enable_vddio
+ gpio6_6_vtrip_sel gpio6_6_ib_mode_sel[1] gpio6_6_ib_mode_sel[0] gpio6_6_out gpio6_6_slew_ctl[1]
+ gpio6_6_slew_ctl[0] gpio6_6_analog_pol gpio6_6_analog_sel gpio6_6_hys_trim gpio6_6_hld_ovr
+ gpio6_6_in_h gpio6_6_enable_h gpio6_6_in gpio6_6_hld_h_n gpio6_6_enable_vdda_h gpio6_6_analog_en
+ gpio6_6_enable_inp_h gpio6_6_enable_vswitch_h gpio6_6_pad_a_noesd_h gpio6_6_pad_a_esd_0_h
+ gpio6_6_pad_a_esd_1_h gpio6_6_zero gpio6_6_one gpio6_7_tie_hi_esd gpio6_7_dm[2]
+ gpio6_7_dm[1] gpio6_7_dm[0] gpio6_7_slow gpio6_7_oe_n gpio6_7_tie_lo_esd gpio6_7_inp_dis
+ gpio6_7_enable_vddio gpio6_7_vtrip_sel gpio6_7_ib_mode_sel[1] gpio6_7_ib_mode_sel[0]
+ gpio6_7_out gpio6_7_slew_ctl[1] gpio6_7_slew_ctl[0] gpio6_7_analog_pol gpio6_7_analog_sel
+ gpio6_7_hys_trim gpio6_7_hld_ovr gpio6_7_in_h gpio6_7_enable_h gpio6_7_in gpio6_7_hld_h_n
+ gpio6_7_enable_vdda_h gpio6_7_analog_en gpio6_7_enable_inp_h gpio6_7_enable_vswitch_h
+ gpio6_7_pad_a_noesd_h gpio6_7_pad_a_esd_0_h gpio6_7_pad_a_esd_1_h gpio6_7_zero gpio6_7_one
+ gpio7_0_tie_lo_esd gpio7_0_in gpio7_0_tie_hi_esd gpio7_0_enable_vddio gpio7_0_slow
+ gpio7_0_pad_a_esd_0_h gpio7_0_pad_a_esd_1_h gpio7_0_pad_a_noesd_h gpio7_0_analog_en
+ gpio7_0_analog_pol gpio7_0_inp_dis gpio7_0_enable_inp_h gpio7_0_enable_h gpio7_0_hld_h_n
+ gpio7_0_analog_sel gpio7_0_dm[2] gpio7_0_dm[1] gpio7_0_dm[0] gpio7_0_hld_ovr gpio7_0_out
+ gpio7_0_enable_vswitch_h gpio7_0_enable_vdda_h gpio7_0_vtrip_sel gpio7_0_ib_mode_sel
+ gpio7_0_oe_n gpio7_0_in_h gpio7_0_zero gpio7_0_one gpio7_1_tie_lo_esd gpio7_1_in
+ gpio7_1_tie_hi_esd gpio7_1_enable_vddio gpio7_1_slow gpio7_1_pad_a_esd_0_h gpio7_1_pad_a_esd_1_h
+ gpio7_1_pad_a_noesd_h gpio7_1_analog_en gpio7_1_analog_pol gpio7_1_inp_dis gpio7_1_enable_inp_h
+ gpio7_1_enable_h gpio7_1_hld_h_n gpio7_1_analog_sel gpio7_1_dm[2] gpio7_1_dm[1]
+ gpio7_1_dm[0] gpio7_1_hld_ovr gpio7_1_out gpio7_1_enable_vswitch_h gpio7_1_enable_vdda_h
+ gpio7_1_vtrip_sel gpio7_1_ib_mode_sel gpio7_1_oe_n gpio7_1_in_h gpio7_1_zero gpio7_1_one
+ gpio7_2_tie_lo_esd gpio7_2_in gpio7_2_tie_hi_esd gpio7_2_enable_vddio gpio7_2_slow
+ gpio7_2_pad_a_esd_0_h gpio7_2_pad_a_esd_1_h gpio7_2_pad_a_noesd_h gpio7_2_analog_en
+ gpio7_2_analog_pol gpio7_2_inp_dis gpio7_2_enable_inp_h gpio7_2_enable_h gpio7_2_hld_h_n
+ gpio7_2_analog_sel gpio7_2_dm[2] gpio7_2_dm[1] gpio7_2_dm[0] gpio7_2_hld_ovr gpio7_2_out
+ gpio7_2_enable_vswitch_h gpio7_2_enable_vdda_h gpio7_2_vtrip_sel gpio7_2_ib_mode_sel
+ gpio7_2_oe_n gpio7_2_in_h gpio7_2_zero gpio7_2_one gpio7_3_tie_lo_esd gpio7_3_in
+ gpio7_3_tie_hi_esd gpio7_3_enable_vddio gpio7_3_slow gpio7_3_pad_a_esd_0_h gpio7_3_pad_a_esd_1_h
+ gpio7_3_pad_a_noesd_h gpio7_3_analog_en gpio7_3_analog_pol gpio7_3_inp_dis gpio7_3_enable_inp_h
+ gpio7_3_enable_h gpio7_3_hld_h_n gpio7_3_analog_sel gpio7_3_dm[2] gpio7_3_dm[1]
+ gpio7_3_dm[0] gpio7_3_hld_ovr gpio7_3_out gpio7_3_enable_vswitch_h gpio7_3_enable_vdda_h
+ gpio7_3_vtrip_sel gpio7_3_ib_mode_sel gpio7_3_oe_n gpio7_3_in_h gpio7_3_zero gpio7_3_one
+ gpio7_4_tie_lo_esd gpio7_4_in gpio7_4_tie_hi_esd gpio7_4_enable_vddio gpio7_4_slow
+ gpio7_4_pad_a_esd_0_h gpio7_4_pad_a_esd_1_h gpio7_4_pad_a_noesd_h gpio7_4_analog_en
+ gpio7_4_analog_pol gpio7_4_inp_dis gpio7_4_enable_inp_h gpio7_4_enable_h gpio7_4_hld_h_n
+ gpio7_4_analog_sel gpio7_4_dm[2] gpio7_4_dm[1] gpio7_4_dm[0] gpio7_4_hld_ovr gpio7_4_out
+ gpio7_4_enable_vswitch_h gpio7_4_enable_vdda_h gpio7_4_vtrip_sel gpio7_4_ib_mode_sel
+ gpio7_4_oe_n gpio7_4_in_h gpio7_4_zero gpio7_4_one gpio7_5_tie_lo_esd gpio7_5_in
+ gpio7_5_tie_hi_esd gpio7_5_enable_vddio gpio7_5_slow gpio7_5_pad_a_esd_0_h gpio7_5_pad_a_esd_1_h
+ gpio7_5_pad_a_noesd_h gpio7_5_analog_en gpio7_5_analog_pol gpio7_5_inp_dis gpio7_5_enable_inp_h
+ gpio7_5_enable_h gpio7_5_hld_h_n gpio7_5_analog_sel gpio7_5_dm[2] gpio7_5_dm[1]
+ gpio7_5_dm[0] gpio7_5_hld_ovr gpio7_5_out gpio7_5_enable_vswitch_h gpio7_5_enable_vdda_h
+ gpio7_5_vtrip_sel gpio7_5_ib_mode_sel gpio7_5_oe_n gpio7_5_in_h gpio7_5_zero gpio7_5_one
+ gpio7_6_tie_lo_esd gpio7_6_in gpio7_6_tie_hi_esd gpio7_6_enable_vddio gpio7_6_slow
+ gpio7_6_pad_a_esd_0_h gpio7_6_pad_a_esd_1_h gpio7_6_pad_a_noesd_h gpio7_6_analog_en
+ gpio7_6_analog_pol gpio7_6_inp_dis gpio7_6_enable_inp_h gpio7_6_enable_h gpio7_6_hld_h_n
+ gpio7_6_analog_sel gpio7_6_dm[2] gpio7_6_dm[1] gpio7_6_dm[0] gpio7_6_hld_ovr gpio7_6_out
+ gpio7_6_enable_vswitch_h gpio7_6_enable_vdda_h gpio7_6_vtrip_sel gpio7_6_ib_mode_sel
+ gpio7_6_oe_n gpio7_6_in_h gpio7_6_zero gpio7_6_one gpio7_7_tie_lo_esd gpio7_7_in
+ gpio7_7_tie_hi_esd gpio7_7_enable_vddio gpio7_7_slow gpio7_7_pad_a_esd_0_h gpio7_7_pad_a_esd_1_h
+ gpio7_7_pad_a_noesd_h gpio7_7_analog_en gpio7_7_analog_pol gpio7_7_inp_dis gpio7_7_enable_inp_h
+ gpio7_7_enable_h gpio7_7_hld_h_n gpio7_7_analog_sel gpio7_7_dm[2] gpio7_7_dm[1]
+ gpio7_7_dm[0] gpio7_7_hld_ovr gpio7_7_out gpio7_7_enable_vswitch_h gpio7_7_enable_vdda_h
+ gpio7_7_vtrip_sel gpio7_7_ib_mode_sel gpio7_7_oe_n gpio7_7_in_h gpio7_7_zero gpio7_7_one
+ muxsplit_sw_hld_vdda_h_n muxsplit_sw_enable_vdda_h muxsplit_sw_switch_aa_sl muxsplit_sw_switch_aa_s0
+ muxsplit_sw_switch_bb_s0 muxsplit_sw_switch_bb_sl muxsplit_sw_switch_bb_sr muxsplit_sw_switch_aa_sr
Xgpio6_3_connects gpio6_3_one gpio6_3_zero gpio6_3_enable_h gpio6_3_tie_hi_esd vcap_w_cpos
+ gpio6_3_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xgpio1_0_pad vcap_w/cneg vddio vssio vssd0 vssa1 vref_w/vddio_q vddio vdda1 vccd0
+ vccd0 gpio1_0 vref_e/amuxbus_a vref_e/amuxbus_b gpio1_0_dm[0] gpio1_0_dm[1] gpio1_0_dm[2]
+ gpio1_0_inp_dis gpio1_0_vtrip_sel gpio1_0_ib_mode_sel[0] gpio1_0_ib_mode_sel[1]
+ gpio1_0_slew_ctl[0] gpio1_0_slew_ctl[1] gpio1_0_hys_trim gpio1_0_hld_ovr gpio1_0_enable_h
+ gpio1_0_hld_h_n gpio1_0_enable_vdda_h gpio1_0_analog_en gpio1_0_enable_inp_h gpio1_0_in
+ gpio1_0_in_h gpio1_0_vinref gpio1_0_out gpio1_0_analog_pol gpio1_0_analog_sel gpio1_0_slow
+ gpio1_0_oe_n gpio1_0_tie_hi_esd gpio1_0_tie_lo_esd gpio1_0_pad_a_esd_0_h gpio1_0_pad_a_esd_1_h
+ gpio1_0_pad_a_noesd_h gpio1_0_enable_vswitch_h gpio1_0_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xgpio3_3_pad gpio3_3_dm[0] gpio3_3_ib_mode_sel gpio3_3_enable_h gpio3_3_enable_inp_h
+ gpio3_3_slow gpio3_3_vtrip_sel gpio3_3_enable_vddio gpio3_3_enable_vdda_h gpio3_3_pad_a_noesd_h
+ gpio3_3_analog_pol gpio3_3_hld_h_n w_572474_1014469# gpio3_3_dm[1] w_575565_1012355#
+ gpio3_3_dm[2] w_572474_1012253# gpio3_3_pad_a_esd_1_h gpio3_3_tie_hi_esd gpio3_3_enable_vswitch_h
+ gpio3_3_tie_lo_esd gpio3_3_oe_n w_575565_1014469# amuxbus_b_n gpio3_3_analog_sel
+ vddio amuxbus_a_n gpio3_3_in_h vddio gpio3_3_inp_dis gpio3_3_out gpio3_3_hld_ovr
+ vccd0 gpio3_3 vccd0 gpio3_3_pad_a_esd_0_h gpio3_3_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio3_3_in vssd0 sky130_ef_io__gpiov2_pad
Xvssio_2_pad vdda1 vssd0 vssa1 vref_e/amuxbus_a vref_e/amuxbus_b vssio_2 vref_w/vddio_q
+ vddio vssio vddio vcap_w/cneg vccd0 vccd0 sky130_ef_io__vssio_hvc_clamped_pad
Xgpio7_6_connects gpio7_6_tie_lo_esd gpio7_6_in gpio7_6_tie_hi_esd gpio7_6_enable_vddio
+ gpio7_6_slow gpio7_6_pad_a_esd_0_h gpio7_6_pad_a_esd_1_h gpio7_6_dm[1] gpio7_6_pad_a_noesd_h
+ gpio7_6_analog_en gpio7_6_dm[0] gpio7_6_analog_pol gpio7_6_inp_dis gpio7_6_enable_inp_h
+ gpio7_6_enable_h gpio7_6_hld_h_n gpio7_6_analog_sel gpio7_6_dm[2] gpio7_6_hld_ovr
+ gpio7_6_out gpio7_6_enable_vswitch_h gpio7_6_enable_vdda_h gpio7_6_vtrip_sel gpio7_6_ib_mode_sel
+ gpio7_6_oe_n gpio7_6_in_h gpio7_6_one gpio7_6_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio5_6_pad gpio5_6_dm[0] gpio5_6_ib_mode_sel gpio5_6_enable_h gpio5_6_enable_inp_h
+ gpio5_6_slow gpio5_6_vtrip_sel gpio5_6_enable_vddio gpio5_6_enable_vdda_h gpio5_6_pad_a_noesd_h
+ gpio5_6_analog_pol gpio5_6_hld_h_n w_21151_791674# gpio5_6_dm[1] w_23367_794765#
+ gpio5_6_dm[2] w_23367_791674# gpio5_6_pad_a_esd_1_h gpio5_6_tie_hi_esd gpio5_6_enable_vswitch_h
+ gpio5_6_tie_lo_esd gpio5_6_oe_n w_21253_794765# vref_w/amuxbus_b gpio5_6_analog_sel
+ vddio vref_w/amuxbus_a gpio5_6_in_h vddio gpio5_6_inp_dis gpio5_6_out gpio5_6_hld_ovr
+ vccd0 gpio5_6 vccd0 gpio5_6_pad_a_esd_0_h gpio5_6_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio5_6_in vssd0 sky130_ef_io__gpiov2_pad
Xvddio_3_pad vdda1 vcap_w/cneg vddio vref_w/vddio_q vssd0 vddio_3 vssa1 vref_e/amuxbus_b
+ vref_e/amuxbus_a vddio vccd0 vssio vccd0 sky130_ef_io__vddio_hvc_clamped_pad
Xgpio0_0_pad gpio0_0_dm[0] gpio0_0_ib_mode_sel gpio0_0_enable_h gpio0_0_enable_inp_h
+ gpio0_0_slow gpio0_0_vtrip_sel gpio0_0_enable_vddio gpio0_0_enable_vdda_h gpio0_0_pad_a_noesd_h
+ gpio0_0_analog_pol gpio0_0_hld_h_n w_694469_78069# gpio0_0_dm[1] w_692355_74752#
+ gpio0_0_dm[2] w_692253_78070# gpio0_0_pad_a_esd_1_h gpio0_0_tie_hi_esd gpio0_0_enable_vswitch_h
+ gpio0_0_tie_lo_esd gpio0_0_oe_n w_694469_74752# vref_e/amuxbus_b gpio0_0_analog_sel
+ vddio vref_e/amuxbus_a gpio0_0_in_h vddio gpio0_0_inp_dis gpio0_0_out gpio0_0_hld_ovr
+ vccd0 gpio0_0 vccd0 gpio0_0_pad_a_esd_0_h gpio0_0_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio0_0_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio2_3_pad gpio2_3_dm[0] gpio2_3_ib_mode_sel gpio2_3_enable_h gpio2_3_enable_inp_h
+ gpio2_3_slow gpio2_3_vtrip_sel gpio2_3_enable_vddio gpio2_3_enable_vdda_h gpio2_3_pad_a_noesd_h
+ gpio2_3_analog_pol gpio2_3_hld_h_n w_694469_825669# gpio2_3_dm[1] w_692355_822352#
+ gpio2_3_dm[2] w_692253_825670# gpio2_3_pad_a_esd_1_h gpio2_3_tie_hi_esd gpio2_3_enable_vswitch_h
+ gpio2_3_tie_lo_esd gpio2_3_oe_n w_694469_822352# vref_e/amuxbus_b gpio2_3_analog_sel
+ vddio vref_e/amuxbus_a gpio2_3_in_h vddio gpio2_3_inp_dis gpio2_3_out gpio2_3_hld_ovr
+ vccd0 gpio2_3 vccd0 gpio2_3_pad_a_esd_0_h gpio2_3_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio2_3_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio4_6_pad gpio4_6_dm[0] gpio4_6_ib_mode_sel gpio4_6_enable_h gpio4_6_enable_inp_h
+ gpio4_6_slow gpio4_6_vtrip_sel gpio4_6_enable_vddio gpio4_6_enable_vdda_h gpio4_6_pad_a_noesd_h
+ gpio4_6_analog_pol gpio4_6_hld_h_n w_101474_1014469# gpio4_6_dm[1] w_104565_1012355#
+ gpio4_6_dm[2] w_101474_1012253# gpio4_6_pad_a_esd_1_h gpio4_6_tie_hi_esd gpio4_6_enable_vswitch_h
+ gpio4_6_tie_lo_esd gpio4_6_oe_n w_104565_1014469# amuxbus_b_n gpio4_6_analog_sel
+ vddio amuxbus_a_n gpio4_6_in_h vddio gpio4_6_inp_dis gpio4_6_out gpio4_6_hld_ovr
+ vccd0 gpio4_6 vccd0 gpio4_6_pad_a_esd_0_h gpio4_6_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio4_6_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio1_1_connects gpio1_1_one gpio1_1_zero gpio1_1_enable_h gpio1_1_tie_hi_esd gpio1_0_vinref
+ gpio1_1_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xvref_w vref_w_ref_sel[4] vref_w_ref_sel[3] vref_w_ref_sel[1] vref_w_vrefgen_en vref_w_hld_h_n
+ vref_w_enable_h vref_w_ref_sel[2] vref_w_ref_sel[0] gpio6_7_vinref vref_w/vddio_q
+ vddio vssio vssa2 vccd0 vccd0 vddio vcap_w/cneg vdda2 vssd0 vref_w/amuxbus_b vref_w/amuxbus_a
+ sky130_fd_io__top_gpiovrefv2
Xvssa2_1_pad vssd0 vssa2 vddio vssa2_1 vddio vssio vccd0 vdda2 vref_w/vddio_q vref_w/amuxbus_a
+ vref_w/amuxbus_b vcap_w/cneg vccd0 sky130_ef_io__vssa_hvc_clamped_pad
Xgpio2_4_connects gpio2_4_tie_lo_esd gpio2_4_in gpio2_4_tie_hi_esd gpio2_4_enable_vddio
+ gpio2_4_slow gpio2_4_pad_a_esd_0_h gpio2_4_pad_a_esd_1_h gpio2_4_dm[1] gpio2_4_pad_a_noesd_h
+ gpio2_4_analog_en gpio2_4_dm[0] gpio2_4_analog_pol gpio2_4_inp_dis gpio2_4_enable_inp_h
+ gpio2_4_enable_h gpio2_4_hld_h_n gpio2_4_analog_sel gpio2_4_dm[2] gpio2_4_hld_ovr
+ gpio2_4_out gpio2_4_enable_vswitch_h gpio2_4_enable_vdda_h gpio2_4_vtrip_sel gpio2_4_ib_mode_sel
+ gpio2_4_oe_n gpio2_4_in_h gpio2_4_one gpio2_4_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio3_7_connects gpio3_7_tie_lo_esd gpio3_7_pad_a_esd_1_h gpio3_7_dm[1] gpio3_7_dm[0]
+ gpio3_7_analog_pol gpio3_7_inp_dis gpio3_7_enable_h gpio3_7_hld_h_n gpio3_7_dm[2]
+ gpio3_7_hld_ovr gpio3_7_out gpio3_7_enable_vswitch_h gpio3_7_enable_vdda_h gpio3_7_vtrip_sel
+ gpio3_7_oe_n gpio3_7_tie_hi_esd gpio3_7_in gpio3_7_enable_vddio gpio3_7_slow gpio3_7_pad_a_esd_0_h
+ gpio3_7_pad_a_noesd_h gpio3_7_analog_en gpio3_7_analog_sel gpio3_7_ib_mode_sel gpio3_7_in_h
+ gpio3_7_zero gpio3_7_one gpio3_7_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio4_0_connects gpio4_0_tie_lo_esd gpio4_0_pad_a_esd_1_h gpio4_0_dm[1] gpio4_0_dm[0]
+ gpio4_0_analog_pol gpio4_0_inp_dis gpio4_0_enable_h gpio4_0_hld_h_n gpio4_0_dm[2]
+ gpio4_0_hld_ovr gpio4_0_out gpio4_0_enable_vswitch_h gpio4_0_enable_vdda_h gpio4_0_vtrip_sel
+ gpio4_0_oe_n gpio4_0_tie_hi_esd gpio4_0_in gpio4_0_enable_vddio gpio4_0_slow gpio4_0_pad_a_esd_0_h
+ gpio4_0_pad_a_noesd_h gpio4_0_analog_en gpio4_0_analog_sel gpio4_0_ib_mode_sel gpio4_0_in_h
+ gpio4_0_zero gpio4_0_one gpio4_0_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio1_3_pad vcap_w/cneg vddio vssio vssd0 vssa1 vref_w/vddio_q vddio vdda1 vccd0
+ vccd0 gpio1_3 vref_e/amuxbus_a vref_e/amuxbus_b gpio1_3_dm[0] gpio1_3_dm[1] gpio1_3_dm[2]
+ gpio1_3_inp_dis gpio1_3_vtrip_sel gpio1_3_ib_mode_sel[0] gpio1_3_ib_mode_sel[1]
+ gpio1_3_slew_ctl[0] gpio1_3_slew_ctl[1] gpio1_3_hys_trim gpio1_3_hld_ovr gpio1_3_enable_h
+ gpio1_3_hld_h_n gpio1_3_enable_vdda_h gpio1_3_analog_en gpio1_3_enable_inp_h gpio1_3_in
+ gpio1_3_in_h gpio1_0_vinref gpio1_3_out gpio1_3_analog_pol gpio1_3_analog_sel gpio1_3_slow
+ gpio1_3_oe_n gpio1_3_tie_hi_esd gpio1_3_tie_lo_esd gpio1_3_pad_a_esd_0_h gpio1_3_pad_a_esd_1_h
+ gpio1_3_pad_a_noesd_h gpio1_3_enable_vswitch_h gpio1_3_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xgpio3_6_pad gpio3_6_dm[0] gpio3_6_ib_mode_sel gpio3_6_enable_h gpio3_6_enable_inp_h
+ gpio3_6_slow gpio3_6_vtrip_sel gpio3_6_enable_vddio gpio3_6_enable_vdda_h gpio3_6_pad_a_noesd_h
+ gpio3_6_analog_pol gpio3_6_hld_h_n w_454474_1014469# gpio3_6_dm[1] w_457565_1012355#
+ gpio3_6_dm[2] w_454474_1012253# gpio3_6_pad_a_esd_1_h gpio3_6_tie_hi_esd gpio3_6_enable_vswitch_h
+ gpio3_6_tie_lo_esd gpio3_6_oe_n w_457565_1014469# amuxbus_b_n gpio3_6_analog_sel
+ vddio amuxbus_a_n gpio3_6_in_h vddio gpio3_6_inp_dis gpio3_6_out gpio3_6_hld_ovr
+ vccd0 gpio3_6 vccd0 gpio3_6_pad_a_esd_0_h gpio3_6_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio3_6_in vssd0 sky130_ef_io__gpiov2_pad
Xvssio_5_pad vdda2 vssd0 vssa2 vref_w/amuxbus_a vref_w/amuxbus_b vssio_5 vref_w/vddio_q
+ vddio vssio vddio vcap_w/cneg vccd0 vccd0 sky130_ef_io__vssio_hvc_clamped_pad
Xgpio5_3_connects gpio5_3_tie_lo_esd gpio5_3_in gpio5_3_tie_hi_esd gpio5_3_enable_vddio
+ gpio5_3_slow gpio5_3_pad_a_esd_0_h gpio5_3_pad_a_esd_1_h gpio5_3_dm[1] gpio5_3_pad_a_noesd_h
+ gpio5_3_analog_en gpio5_3_dm[0] gpio5_3_analog_pol gpio5_3_inp_dis gpio5_3_enable_inp_h
+ gpio5_3_enable_h gpio5_3_hld_h_n gpio5_3_analog_sel gpio5_3_dm[2] gpio5_3_hld_ovr
+ gpio5_3_out gpio5_3_enable_vswitch_h gpio5_3_enable_vdda_h gpio5_3_vtrip_sel gpio5_3_ib_mode_sel
+ gpio5_3_oe_n gpio5_3_in_h gpio5_3_one gpio5_3_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xmuxsplit_se sio_amuxbus_a vref_e/amuxbus_a sio_amuxbus_b vref_e/amuxbus_b muxsplit_se_enable_vdda_h
+ muxsplit_se_hld_vdda_h_n muxsplit_se_switch_aa_s0 muxsplit_se_switch_aa_sl muxsplit_se_switch_aa_sr
+ muxsplit_se_switch_bb_s0 muxsplit_se_switch_bb_sl muxsplit_se_switch_bb_sr vssd0
+ vssio vddio vccd0 vref_w/vddio_q vddio vccd0 w_707299_42182# w_700999_42182# vdda3
+ vssa3 vcap_w/cneg sky130_fd_io__top_amuxsplitv2
Xvssa1_1_pad vssd0 vssa1 vddio vssa1_1 vddio vssio vccd0 vdda1 vref_w/vddio_q vref_e/amuxbus_a
+ vref_e/amuxbus_b vcap_w/cneg vccd0 sky130_ef_io__vssa_hvc_clamped_pad
Xgpio6_6_connects gpio6_6_one gpio6_6_zero gpio6_6_enable_h gpio6_6_tie_hi_esd gpio6_7_vinref
+ gpio6_6_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xvddio_6_pad vdda2 vcap_w/cneg vddio vref_w/vddio_q vssd0 vddio_6 vssa2 vref_w/amuxbus_b
+ vref_w/amuxbus_a vddio vccd0 vssio vccd0 sky130_ef_io__vddio_hvc_clamped_pad
Xgpio0_3_pad gpio0_3_dm[0] gpio0_3_ib_mode_sel gpio0_3_enable_h gpio0_3_enable_inp_h
+ gpio0_3_slow gpio0_3_vtrip_sel gpio0_3_enable_vddio gpio0_3_enable_vdda_h gpio0_3_pad_a_noesd_h
+ gpio0_3_analog_pol gpio0_3_hld_h_n w_694469_141069# gpio0_3_dm[1] w_692355_137752#
+ gpio0_3_dm[2] w_692253_141070# gpio0_3_pad_a_esd_1_h gpio0_3_tie_hi_esd gpio0_3_enable_vswitch_h
+ gpio0_3_tie_lo_esd gpio0_3_oe_n w_694469_137752# vref_e/amuxbus_b gpio0_3_analog_sel
+ vddio vref_e/amuxbus_a gpio0_3_in_h vddio gpio0_3_inp_dis gpio0_3_out gpio0_3_hld_ovr
+ vccd0 gpio0_3 vccd0 gpio0_3_pad_a_esd_0_h gpio0_3_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio0_3_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio8_2_connects gpio8_2_tie_lo_esd gpio8_2_pad_a_esd_1_h gpio8_2_dm[1] gpio8_2_dm[0]
+ gpio8_2_analog_pol gpio8_2_inp_dis gpio8_2_enable_h gpio8_2_hld_h_n gpio8_2_dm[2]
+ gpio8_2_hld_ovr gpio8_2_out gpio8_2_enable_vswitch_h gpio8_2_enable_vdda_h gpio8_2_vtrip_sel
+ gpio8_2_oe_n gpio8_2_tie_hi_esd gpio8_2_in gpio8_2_enable_vddio gpio8_2_slow gpio8_2_pad_a_esd_0_h
+ gpio8_2_pad_a_noesd_h gpio8_2_analog_en gpio8_2_analog_sel gpio8_2_ib_mode_sel gpio8_2_in_h
+ gpio8_2_zero gpio8_2_one gpio8_2_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio2_6_pad gpio2_6_dm[0] gpio2_6_ib_mode_sel gpio2_6_enable_h gpio2_6_enable_inp_h
+ gpio2_6_slow gpio2_6_vtrip_sel gpio2_6_enable_vddio gpio2_6_enable_vdda_h gpio2_6_pad_a_noesd_h
+ gpio2_6_analog_pol gpio2_6_hld_h_n w_694469_908669# gpio2_6_dm[1] w_692355_905352#
+ gpio2_6_dm[2] w_692253_908670# gpio2_6_pad_a_esd_1_h gpio2_6_tie_hi_esd gpio2_6_enable_vswitch_h
+ gpio2_6_tie_lo_esd gpio2_6_oe_n w_694469_905352# vref_e/amuxbus_b gpio2_6_analog_sel
+ vddio vref_e/amuxbus_a gpio2_6_in_h vddio gpio2_6_inp_dis gpio2_6_out gpio2_6_hld_ovr
+ vccd0 gpio2_6 vccd0 gpio2_6_pad_a_esd_0_h gpio2_6_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio2_6_in vssd0 sky130_ef_io__gpiov2_pad
Xxo0_pad vccd0 vref_w/vddio_q vccd0 vcap_w/cneg vssd0 sio_amuxbus_b sio_amuxbus_a
+ xo0_core vssa3 vddio vddio vdda3 vssio xo0 sky130_fd_io__top_analog_pad
Xgpio8_2_pad gpio8_2_dm[0] gpio8_2_ib_mode_sel gpio8_2_enable_h gpio8_2_enable_inp_h
+ gpio8_2_slow gpio8_2_vtrip_sel gpio8_2_enable_vddio gpio8_2_enable_vdda_h gpio8_2_pad_a_noesd_h
+ gpio8_2_analog_pol gpio8_2_hld_h_n w_163469_21253# gpio8_2_dm[1] w_160152_23367#
+ gpio8_2_dm[2] w_163469_23367# gpio8_2_pad_a_esd_1_h gpio8_2_tie_hi_esd gpio8_2_enable_vswitch_h
+ gpio8_2_tie_lo_esd gpio8_2_oe_n w_160152_21253# sio_amuxbus_b gpio8_2_analog_sel
+ vddio sio_amuxbus_a gpio8_2_in_h vddio gpio8_2_inp_dis gpio8_2_out gpio8_2_hld_ovr
+ vccd0 gpio8_2 vccd0 gpio8_2_pad_a_esd_0_h gpio8_2_analog_en vssio vdda3 vref_w/vddio_q
+ vcap_w/cneg vssa3 gpio8_2_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio0_1_connects gpio0_1_tie_lo_esd gpio0_1_in gpio0_1_tie_hi_esd gpio0_1_enable_vddio
+ gpio0_1_slow gpio0_1_pad_a_esd_0_h gpio0_1_pad_a_esd_1_h gpio0_1_dm[1] gpio0_1_pad_a_noesd_h
+ gpio0_1_analog_en gpio0_1_dm[0] gpio0_1_analog_pol gpio0_1_inp_dis gpio0_1_enable_inp_h
+ gpio0_1_enable_h gpio0_1_hld_h_n gpio0_1_analog_sel gpio0_1_dm[2] gpio0_1_hld_ovr
+ gpio0_1_out gpio0_1_enable_vswitch_h gpio0_1_enable_vdda_h gpio0_1_vtrip_sel gpio0_1_ib_mode_sel
+ gpio0_1_oe_n gpio0_1_in_h gpio0_1_one gpio0_1_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio1_4_connects gpio1_4_one gpio1_4_zero gpio1_4_enable_h gpio1_4_tie_hi_esd vcap_e_cpos
+ gpio1_4_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xgpio1_6_pad vcap_w/cneg vddio vssio vssd0 vssa1 vref_w/vddio_q vddio vdda1 vccd0
+ vccd0 gpio1_6 vref_e/amuxbus_a vref_e/amuxbus_b gpio1_6_dm[0] gpio1_6_dm[1] gpio1_6_dm[2]
+ gpio1_6_inp_dis gpio1_6_vtrip_sel gpio1_6_ib_mode_sel[0] gpio1_6_ib_mode_sel[1]
+ gpio1_6_slew_ctl[0] gpio1_6_slew_ctl[1] gpio1_6_hys_trim gpio1_6_hld_ovr gpio1_6_enable_h
+ gpio1_6_hld_h_n gpio1_6_enable_vdda_h gpio1_6_analog_en gpio1_6_enable_inp_h gpio1_6_in
+ gpio1_6_in_h vcap_e_cpos gpio1_6_out gpio1_6_analog_pol gpio1_6_analog_sel gpio1_6_slow
+ gpio1_6_oe_n gpio1_6_tie_hi_esd gpio1_6_tie_lo_esd gpio1_6_pad_a_esd_0_h gpio1_6_pad_a_esd_1_h
+ gpio1_6_pad_a_noesd_h gpio1_6_enable_vswitch_h gpio1_6_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xgpio2_7_connects gpio2_7_tie_lo_esd gpio2_7_in gpio2_7_tie_hi_esd gpio2_7_enable_vddio
+ gpio2_7_slow gpio2_7_pad_a_esd_0_h gpio2_7_pad_a_esd_1_h gpio2_7_dm[1] gpio2_7_pad_a_noesd_h
+ gpio2_7_analog_en gpio2_7_dm[0] gpio2_7_analog_pol gpio2_7_inp_dis gpio2_7_enable_inp_h
+ gpio2_7_enable_h gpio2_7_hld_h_n gpio2_7_analog_sel gpio2_7_dm[2] gpio2_7_hld_ovr
+ gpio2_7_out gpio2_7_enable_vswitch_h gpio2_7_enable_vdda_h gpio2_7_vtrip_sel gpio2_7_ib_mode_sel
+ gpio2_7_oe_n gpio2_7_in_h gpio2_7_one gpio2_7_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xvssio_8_pad vdda3 vssd0 vssa3 sio_amuxbus_a sio_amuxbus_b vssio_8 vref_w/vddio_q
+ vddio vssio vddio vcap_w/cneg vccd0 vccd0 sky130_ef_io__vssio_hvc_clamped_pad
Xgpio3_0_connects gpio3_0_tie_lo_esd gpio3_0_pad_a_esd_1_h gpio3_0_dm[1] gpio3_0_dm[0]
+ gpio3_0_analog_pol gpio3_0_inp_dis gpio3_0_enable_h gpio3_0_hld_h_n gpio3_0_dm[2]
+ gpio3_0_hld_ovr gpio3_0_out gpio3_0_enable_vswitch_h gpio3_0_enable_vdda_h gpio3_0_vtrip_sel
+ gpio3_0_oe_n gpio3_0_tie_hi_esd gpio3_0_in gpio3_0_enable_vddio gpio3_0_slow gpio3_0_pad_a_esd_0_h
+ gpio3_0_pad_a_noesd_h gpio3_0_analog_en gpio3_0_analog_sel gpio3_0_ib_mode_sel gpio3_0_in_h
+ gpio3_0_zero gpio3_0_one gpio3_0_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xvccd2_2_pad vdda2 vccd0 vssd2[5] vddio vref_w/amuxbus_b vddio vssio vref_w/amuxbus_a
+ vccd0 vccd2_2 vccd2[5] vssd0 vssa2 vref_w/vddio_q vcap_w/cneg sky130_ef_io__vccd_lvc_clamped3_pad
Xgpio7_2_pad gpio7_2_dm[0] gpio7_2_ib_mode_sel gpio7_2_enable_h gpio7_2_enable_inp_h
+ gpio7_2_slow gpio7_2_vtrip_sel gpio7_2_enable_vddio gpio7_2_enable_vdda_h gpio7_2_pad_a_noesd_h
+ gpio7_2_analog_pol gpio7_2_hld_h_n w_21151_233074# gpio7_2_dm[1] w_23367_236165#
+ gpio7_2_dm[2] w_23367_233074# gpio7_2_pad_a_esd_1_h gpio7_2_tie_hi_esd gpio7_2_enable_vswitch_h
+ gpio7_2_tie_lo_esd gpio7_2_oe_n w_21253_236165# vref_w/amuxbus_b gpio7_2_analog_sel
+ vddio vref_w/amuxbus_a gpio7_2_in_h vddio gpio7_2_inp_dis gpio7_2_out gpio7_2_hld_ovr
+ vccd0 gpio7_2 vccd0 gpio7_2_pad_a_esd_0_h gpio7_2_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio7_2_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio4_3_connects gpio4_3_tie_lo_esd gpio4_3_pad_a_esd_1_h gpio4_3_dm[1] gpio4_3_dm[0]
+ gpio4_3_analog_pol gpio4_3_inp_dis gpio4_3_enable_h gpio4_3_hld_h_n gpio4_3_dm[2]
+ gpio4_3_hld_ovr gpio4_3_out gpio4_3_enable_vswitch_h gpio4_3_enable_vdda_h gpio4_3_vtrip_sel
+ gpio4_3_oe_n gpio4_3_tie_hi_esd gpio4_3_in gpio4_3_enable_vddio gpio4_3_slow gpio4_3_pad_a_esd_0_h
+ gpio4_3_pad_a_noesd_h gpio4_3_analog_en gpio4_3_analog_sel gpio4_3_ib_mode_sel gpio4_3_in_h
+ gpio4_3_zero gpio4_3_one gpio4_3_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xvddio_9_pad vdda3 vcap_w/cneg vddio vref_w/vddio_q vssd0 vddio_9 vssa3 sio_amuxbus_b
+ sio_amuxbus_a vddio vccd0 vssio vccd0 sky130_ef_io__vddio_hvc_clamped_pad
Xgpio5_6_connects gpio5_6_tie_lo_esd gpio5_6_in gpio5_6_tie_hi_esd gpio5_6_enable_vddio
+ gpio5_6_slow gpio5_6_pad_a_esd_0_h gpio5_6_pad_a_esd_1_h gpio5_6_dm[1] gpio5_6_pad_a_noesd_h
+ gpio5_6_analog_en gpio5_6_dm[0] gpio5_6_analog_pol gpio5_6_inp_dis gpio5_6_enable_inp_h
+ gpio5_6_enable_h gpio5_6_hld_h_n gpio5_6_analog_sel gpio5_6_dm[2] gpio5_6_hld_ovr
+ gpio5_6_out gpio5_6_enable_vswitch_h gpio5_6_enable_vdda_h gpio5_6_vtrip_sel gpio5_6_ib_mode_sel
+ gpio5_6_oe_n gpio5_6_in_h gpio5_6_one gpio5_6_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio0_6_pad gpio0_6_dm[0] gpio0_6_ib_mode_sel gpio0_6_enable_h gpio0_6_enable_inp_h
+ gpio0_6_slow gpio0_6_vtrip_sel gpio0_6_enable_vddio gpio0_6_enable_vdda_h gpio0_6_pad_a_noesd_h
+ gpio0_6_analog_pol gpio0_6_hld_h_n w_694469_244069# gpio0_6_dm[1] w_692355_240752#
+ gpio0_6_dm[2] w_692253_244070# gpio0_6_pad_a_esd_1_h gpio0_6_tie_hi_esd gpio0_6_enable_vswitch_h
+ gpio0_6_tie_lo_esd gpio0_6_oe_n w_694469_240752# vref_e/amuxbus_b gpio0_6_analog_sel
+ vddio vref_e/amuxbus_a gpio0_6_in_h vddio gpio0_6_inp_dis gpio0_6_out gpio0_6_hld_ovr
+ vccd0 gpio0_6 vccd0 gpio0_6_pad_a_esd_0_h gpio0_6_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio0_6_in vssd0 sky130_ef_io__gpiov2_pad
Xvccd1_2_pad vdda0 vccd0 vssd1[5] vddio amuxbus_b_n vddio vssio amuxbus_a_n vccd0
+ vccd1_2 vccd1[5] vssd0 vssa0 vref_w/vddio_q vcap_w/cneg sky130_ef_io__vccd_lvc_clamped3_pad
Xgpio7_2_connects gpio7_2_tie_lo_esd gpio7_2_in gpio7_2_tie_hi_esd gpio7_2_enable_vddio
+ gpio7_2_slow gpio7_2_pad_a_esd_0_h gpio7_2_pad_a_esd_1_h gpio7_2_dm[1] gpio7_2_pad_a_noesd_h
+ gpio7_2_analog_en gpio7_2_dm[0] gpio7_2_analog_pol gpio7_2_inp_dis gpio7_2_enable_inp_h
+ gpio7_2_enable_h gpio7_2_hld_h_n gpio7_2_analog_sel gpio7_2_dm[2] gpio7_2_hld_ovr
+ gpio7_2_out gpio7_2_enable_vswitch_h gpio7_2_enable_vdda_h gpio7_2_vtrip_sel gpio7_2_ib_mode_sel
+ gpio7_2_oe_n gpio7_2_in_h gpio7_2_one gpio7_2_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio6_2_pad vcap_w/cneg vddio vssio vssd0 vssa2 vref_w/vddio_q vddio vdda2 vccd0
+ vccd0 gpio6_2 vref_w/amuxbus_a vref_w/amuxbus_b gpio6_2_dm[0] gpio6_2_dm[1] gpio6_2_dm[2]
+ gpio6_2_inp_dis gpio6_2_vtrip_sel gpio6_2_ib_mode_sel[0] gpio6_2_ib_mode_sel[1]
+ gpio6_2_slew_ctl[0] gpio6_2_slew_ctl[1] gpio6_2_hys_trim gpio6_2_hld_ovr gpio6_2_enable_h
+ gpio6_2_hld_h_n gpio6_2_enable_vdda_h gpio6_2_analog_en gpio6_2_enable_inp_h gpio6_2_in
+ gpio6_2_in_h vcap_w_cpos gpio6_2_out gpio6_2_analog_pol gpio6_2_analog_sel gpio6_2_slow
+ gpio6_2_oe_n gpio6_2_tie_hi_esd gpio6_2_tie_lo_esd gpio6_2_pad_a_esd_0_h gpio6_2_pad_a_esd_1_h
+ gpio6_2_pad_a_noesd_h gpio6_2_enable_vswitch_h gpio6_2_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xgpio8_5_pad gpio8_5_dm[0] gpio8_5_ib_mode_sel gpio8_5_enable_h gpio8_5_enable_inp_h
+ gpio8_5_slow gpio8_5_vtrip_sel gpio8_5_enable_vddio gpio8_5_enable_vdda_h gpio8_5_pad_a_noesd_h
+ gpio8_5_analog_pol gpio8_5_hld_h_n w_412469_21253# gpio8_5_dm[1] w_409152_23367#
+ gpio8_5_dm[2] w_412469_23367# gpio8_5_pad_a_esd_1_h gpio8_5_tie_hi_esd gpio8_5_enable_vswitch_h
+ gpio8_5_tie_lo_esd gpio8_5_oe_n w_409152_21253# sio_amuxbus_b gpio8_5_analog_sel
+ vddio sio_amuxbus_a gpio8_5_in_h vddio gpio8_5_inp_dis gpio8_5_out gpio8_5_hld_ovr
+ vccd0 gpio8_5 vccd0 gpio8_5_pad_a_esd_0_h gpio8_5_analog_en vssio vdda3 vref_w/vddio_q
+ vcap_w/cneg vssa3 gpio8_5_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio8_5_connects gpio8_5_tie_lo_esd gpio8_5_pad_a_esd_1_h gpio8_5_dm[1] gpio8_5_dm[0]
+ gpio8_5_analog_pol gpio8_5_inp_dis gpio8_5_enable_h gpio8_5_hld_h_n gpio8_5_dm[2]
+ gpio8_5_hld_ovr gpio8_5_out gpio8_5_enable_vswitch_h gpio8_5_enable_vdda_h gpio8_5_vtrip_sel
+ gpio8_5_oe_n gpio8_5_tie_hi_esd gpio8_5_in gpio8_5_enable_vddio gpio8_5_slow gpio8_5_pad_a_esd_0_h
+ gpio8_5_pad_a_noesd_h gpio8_5_analog_en gpio8_5_analog_sel gpio8_5_ib_mode_sel gpio8_5_in_h
+ gpio8_5_zero gpio8_5_one gpio8_5_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xmuxsplit_ne vref_e/amuxbus_a amuxbus_a_n vref_e/amuxbus_b amuxbus_b_n muxsplit_ne_enable_vdda_h
+ muxsplit_ne_hld_vdda_h_n muxsplit_ne_switch_aa_s0 muxsplit_ne_switch_aa_sl muxsplit_ne_switch_aa_sr
+ muxsplit_ne_switch_bb_s0 muxsplit_ne_switch_bb_sl muxsplit_ne_switch_bb_sr vssd0
+ vssio vddio vccd0 vref_w/vddio_q vddio vccd0 w_707299_989382# w_700999_989382# vdda0
+ vssa0 vcap_w/cneg sky130_fd_io__top_amuxsplitv2
Xgpio5_2_pad gpio5_2_dm[0] gpio5_2_ib_mode_sel gpio5_2_enable_h gpio5_2_enable_inp_h
+ gpio5_2_slow gpio5_2_vtrip_sel gpio5_2_enable_vddio gpio5_2_enable_vdda_h gpio5_2_pad_a_noesd_h
+ gpio5_2_analog_pol gpio5_2_hld_h_n w_21151_895674# gpio5_2_dm[1] w_23367_898765#
+ gpio5_2_dm[2] w_23367_895674# gpio5_2_pad_a_esd_1_h gpio5_2_tie_hi_esd gpio5_2_enable_vswitch_h
+ gpio5_2_tie_lo_esd gpio5_2_oe_n w_21253_898765# vref_w/amuxbus_b gpio5_2_analog_sel
+ vddio vref_w/amuxbus_a gpio5_2_in_h vddio gpio5_2_inp_dis gpio5_2_out gpio5_2_hld_ovr
+ vccd0 gpio5_2 vccd0 gpio5_2_pad_a_esd_0_h gpio5_2_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio5_2_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio0_4_connects gpio0_4_tie_lo_esd gpio0_4_in gpio0_4_tie_hi_esd gpio0_4_enable_vddio
+ gpio0_4_slow gpio0_4_pad_a_esd_0_h gpio0_4_pad_a_esd_1_h gpio0_4_dm[1] gpio0_4_pad_a_noesd_h
+ gpio0_4_analog_en gpio0_4_dm[0] gpio0_4_analog_pol gpio0_4_inp_dis gpio0_4_enable_inp_h
+ gpio0_4_enable_h gpio0_4_hld_h_n gpio0_4_analog_sel gpio0_4_dm[2] gpio0_4_hld_ovr
+ gpio0_4_out gpio0_4_enable_vswitch_h gpio0_4_enable_vdda_h gpio0_4_vtrip_sel gpio0_4_ib_mode_sel
+ gpio0_4_oe_n gpio0_4_in_h gpio0_4_one gpio0_4_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio7_5_pad gpio7_5_dm[0] gpio7_5_ib_mode_sel gpio7_5_enable_h gpio7_5_enable_inp_h
+ gpio7_5_slow gpio7_5_vtrip_sel gpio7_5_enable_vddio gpio7_5_enable_vdda_h gpio7_5_pad_a_noesd_h
+ gpio7_5_analog_pol gpio7_5_hld_h_n w_21151_127074# gpio7_5_dm[1] w_23367_130165#
+ gpio7_5_dm[2] w_23367_127074# gpio7_5_pad_a_esd_1_h gpio7_5_tie_hi_esd gpio7_5_enable_vswitch_h
+ gpio7_5_tie_lo_esd gpio7_5_oe_n w_21253_130165# vref_w/amuxbus_b gpio7_5_analog_sel
+ vddio vref_w/amuxbus_a gpio7_5_in_h vddio gpio7_5_inp_dis gpio7_5_out gpio7_5_hld_ovr
+ vccd0 gpio7_5 vccd0 gpio7_5_pad_a_esd_0_h gpio7_5_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio7_5_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio1_7_connects gpio1_7_one gpio1_7_zero gpio1_7_enable_h gpio1_7_tie_hi_esd vcap_e_cpos
+ gpio1_7_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xgpio2_0_connects gpio2_0_tie_lo_esd gpio2_0_in gpio2_0_tie_hi_esd gpio2_0_enable_vddio
+ gpio2_0_slow gpio2_0_pad_a_esd_0_h gpio2_0_pad_a_esd_1_h gpio2_0_dm[1] gpio2_0_pad_a_noesd_h
+ gpio2_0_analog_en gpio2_0_dm[0] gpio2_0_analog_pol gpio2_0_inp_dis gpio2_0_enable_inp_h
+ gpio2_0_enable_h gpio2_0_hld_h_n gpio2_0_analog_sel gpio2_0_dm[2] gpio2_0_hld_ovr
+ gpio2_0_out gpio2_0_enable_vswitch_h gpio2_0_enable_vdda_h gpio2_0_vtrip_sel gpio2_0_ib_mode_sel
+ gpio2_0_oe_n gpio2_0_in_h gpio2_0_one gpio2_0_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio3_3_connects gpio3_3_tie_lo_esd gpio3_3_pad_a_esd_1_h gpio3_3_dm[1] gpio3_3_dm[0]
+ gpio3_3_analog_pol gpio3_3_inp_dis gpio3_3_enable_h gpio3_3_hld_h_n gpio3_3_dm[2]
+ gpio3_3_hld_ovr gpio3_3_out gpio3_3_enable_vswitch_h gpio3_3_enable_vdda_h gpio3_3_vtrip_sel
+ gpio3_3_oe_n gpio3_3_tie_hi_esd gpio3_3_in gpio3_3_enable_vddio gpio3_3_slow gpio3_3_pad_a_esd_0_h
+ gpio3_3_pad_a_noesd_h gpio3_3_analog_en gpio3_3_analog_sel gpio3_3_ib_mode_sel gpio3_3_in_h
+ gpio3_3_zero gpio3_3_one gpio3_3_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xanalog_0_pad vccd0 vref_w/vddio_q vccd0 vcap_w/cneg vssd0 amuxbus_b_n amuxbus_a_n
+ analog_0_core vssa0 vddio vddio vdda0 vssio analog_0 sky130_fd_io__top_analog_pad
Xgpio4_2_pad gpio4_2_dm[0] gpio4_2_ib_mode_sel gpio4_2_enable_h gpio4_2_enable_inp_h
+ gpio4_2_slow gpio4_2_vtrip_sel gpio4_2_enable_vddio gpio4_2_enable_vdda_h gpio4_2_pad_a_noesd_h
+ gpio4_2_analog_pol gpio4_2_hld_h_n w_243474_1014469# gpio4_2_dm[1] w_246565_1012355#
+ gpio4_2_dm[2] w_243474_1012253# gpio4_2_pad_a_esd_1_h gpio4_2_tie_hi_esd gpio4_2_enable_vswitch_h
+ gpio4_2_tie_lo_esd gpio4_2_oe_n w_246565_1014469# amuxbus_b_n gpio4_2_analog_sel
+ vddio amuxbus_a_n gpio4_2_in_h vddio gpio4_2_inp_dis gpio4_2_out gpio4_2_hld_ovr
+ vccd0 gpio4_2 vccd0 gpio4_2_pad_a_esd_0_h gpio4_2_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio4_2_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio4_6_connects gpio4_6_tie_lo_esd gpio4_6_pad_a_esd_1_h gpio4_6_dm[1] gpio4_6_dm[0]
+ gpio4_6_analog_pol gpio4_6_inp_dis gpio4_6_enable_h gpio4_6_hld_h_n gpio4_6_dm[2]
+ gpio4_6_hld_ovr gpio4_6_out gpio4_6_enable_vswitch_h gpio4_6_enable_vdda_h gpio4_6_vtrip_sel
+ gpio4_6_oe_n gpio4_6_tie_hi_esd gpio4_6_in gpio4_6_enable_vddio gpio4_6_slow gpio4_6_pad_a_esd_0_h
+ gpio4_6_pad_a_noesd_h gpio4_6_analog_en gpio4_6_analog_sel gpio4_6_ib_mode_sel gpio4_6_in_h
+ gpio4_6_zero gpio4_6_one gpio4_6_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio6_5_pad vcap_w/cneg vddio vssio vssd0 vssa2 vref_w/vddio_q vddio vdda2 vccd0
+ vccd0 gpio6_5 vref_w/amuxbus_a vref_w/amuxbus_b gpio6_5_dm[0] gpio6_5_dm[1] gpio6_5_dm[2]
+ gpio6_5_inp_dis gpio6_5_vtrip_sel gpio6_5_ib_mode_sel[0] gpio6_5_ib_mode_sel[1]
+ gpio6_5_slew_ctl[0] gpio6_5_slew_ctl[1] gpio6_5_hys_trim gpio6_5_hld_ovr gpio6_5_enable_h
+ gpio6_5_hld_h_n gpio6_5_enable_vdda_h gpio6_5_analog_en gpio6_5_enable_inp_h gpio6_5_in
+ gpio6_5_in_h gpio6_7_vinref gpio6_5_out gpio6_5_analog_pol gpio6_5_analog_sel gpio6_5_slow
+ gpio6_5_oe_n gpio6_5_tie_hi_esd gpio6_5_tie_lo_esd gpio6_5_pad_a_esd_0_h gpio6_5_pad_a_esd_1_h
+ gpio6_5_pad_a_noesd_h gpio6_5_enable_vswitch_h gpio6_5_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xvssd2_2_pad vdda2 vcap_w/cneg vssd2[4] vccd0 vssd0 vssa2 vref_w/amuxbus_b vref_w/amuxbus_a
+ vssd2_2 vddio vddio vccd0 vref_w/vddio_q vssio vccd2[4] sky130_ef_io__vssd_lvc_clamped3_pad
Xsio_macro_pads vssa3 vddio vccd0 vccd0 vdda3 vref_w/vddio_q vssd0 vssio vddio vcap_w/cneg
+ sio0 sio1 sio_amuxbus_b sio_amuxbus_a sio_vreg_en_refgen sio_hld_h_n_refgen sio_voh_sel[0]
+ sio_voh_sel[1] sio_voh_sel[2] sio_vohref sio_enable_vdda_h sio_vtrip_sel_refgen
+ sio_dft_refgen sio_dm1[1] sio_dm1[2] sio_dm1[0] sio_dm0[0] sio_dm0[1] sio_dm0[2]
+ sio_voutref_dft sio_ibuf_sel_refgen sio_vref_sel[0] sio_pad_a_esd_1_h[0] sio_ibuf_sel[1]
+ sio_vinref_dft sio_pad_a_esd_1_h[1] sio_pad_a_esd_0_h[1] sio_vref_sel[1] sio_pad_a_esd_0_h[0]
+ sio_pad_a_noesd_h[0] sio_pad_a_noesd_h[1] sio_inp_dis[1] sio_inp_dis[0] sio_tie_lo_esd[0]
+ sio_tie_lo_esd[1] sio_out[1] sio_out[0] sio_vtrip_sel[0] sio_vtrip_sel[1] sio_enable_h
+ sio_vreg_en[0] sio_vreg_en[1] sio_slow[1] sio_slow[0] sio_oe_n[0] sio_oe_n[1] sio_in_h[1]
+ sio_in_h[0] sio_in[0] sio_in[1] sio_hld_ovr[1] sio_hld_ovr[0] sio_hld_h_n[1] sio_hld_h_n[0]
+ sio_ibuf_sel[0] sky130_fd_io__top_sio_macro
Xgpio6_2_connects gpio6_2_one gpio6_2_zero gpio6_2_enable_h gpio6_2_tie_hi_esd vcap_w_cpos
+ gpio6_2_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xgpio7_5_connects gpio7_5_tie_lo_esd gpio7_5_in gpio7_5_tie_hi_esd gpio7_5_enable_vddio
+ gpio7_5_slow gpio7_5_pad_a_esd_0_h gpio7_5_pad_a_esd_1_h gpio7_5_dm[1] gpio7_5_pad_a_noesd_h
+ gpio7_5_analog_en gpio7_5_dm[0] gpio7_5_analog_pol gpio7_5_inp_dis gpio7_5_enable_inp_h
+ gpio7_5_enable_h gpio7_5_hld_h_n gpio7_5_analog_sel gpio7_5_dm[2] gpio7_5_hld_ovr
+ gpio7_5_out gpio7_5_enable_vswitch_h gpio7_5_enable_vdda_h gpio7_5_vtrip_sel gpio7_5_ib_mode_sel
+ gpio7_5_oe_n gpio7_5_in_h gpio7_5_one gpio7_5_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio3_2_pad gpio3_2_dm[0] gpio3_2_ib_mode_sel gpio3_2_enable_h gpio3_2_enable_inp_h
+ gpio3_2_slow gpio3_2_vtrip_sel gpio3_2_enable_vddio gpio3_2_enable_vdda_h gpio3_2_pad_a_noesd_h
+ gpio3_2_analog_pol gpio3_2_hld_h_n w_596474_1014469# gpio3_2_dm[1] w_599565_1012355#
+ gpio3_2_dm[2] w_596474_1012253# gpio3_2_pad_a_esd_1_h gpio3_2_tie_hi_esd gpio3_2_enable_vswitch_h
+ gpio3_2_tie_lo_esd gpio3_2_oe_n w_599565_1014469# amuxbus_b_n gpio3_2_analog_sel
+ vddio amuxbus_a_n gpio3_2_in_h vddio gpio3_2_inp_dis gpio3_2_out gpio3_2_hld_ovr
+ vccd0 gpio3_2 vccd0 gpio3_2_pad_a_esd_0_h gpio3_2_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio3_2_in vssd0 sky130_ef_io__gpiov2_pad
Xvssio_1_pad vdda1 vssd0 vssa1 vref_e/amuxbus_a vref_e/amuxbus_b vssio_1 vref_w/vddio_q
+ vddio vssio vddio vcap_w/cneg vccd0 vccd0 sky130_ef_io__vssio_hvc_clamped_pad
Xvssd1_2_pad vdda0 vcap_w/cneg vssd1[4] vccd0 vssd0 vssa0 amuxbus_b_n amuxbus_a_n
+ vssd1_2 vddio vddio vccd0 vref_w/vddio_q vssio vccd1[4] sky130_ef_io__vssd_lvc_clamped3_pad
Xgpio5_5_pad gpio5_5_dm[0] gpio5_5_ib_mode_sel gpio5_5_enable_h gpio5_5_enable_inp_h
+ gpio5_5_slow gpio5_5_vtrip_sel gpio5_5_enable_vddio gpio5_5_enable_vdda_h gpio5_5_pad_a_noesd_h
+ gpio5_5_analog_pol gpio5_5_hld_h_n w_21151_812674# gpio5_5_dm[1] w_23367_815765#
+ gpio5_5_dm[2] w_23367_812674# gpio5_5_pad_a_esd_1_h gpio5_5_tie_hi_esd gpio5_5_enable_vswitch_h
+ gpio5_5_tie_lo_esd gpio5_5_oe_n w_21253_815765# vref_w/amuxbus_b gpio5_5_analog_sel
+ vddio vref_w/amuxbus_a gpio5_5_in_h vddio gpio5_5_inp_dis gpio5_5_out gpio5_5_hld_ovr
+ vccd0 gpio5_5 vccd0 gpio5_5_pad_a_esd_0_h gpio5_5_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio5_5_in vssd0 sky130_ef_io__gpiov2_pad
Xvssa3_0_pad vssd0 vssa3 vddio vssa3_0 vddio vssio vccd0 vdda3 vref_w/vddio_q sio_amuxbus_a
+ sio_amuxbus_b vcap_w/cneg vccd0 sky130_ef_io__vssa_hvc_clamped_pad
Xvddio_2_pad vdda1 vcap_w/cneg vddio vref_w/vddio_q vssd0 vddio_2 vssa1 vref_e/amuxbus_b
+ vref_e/amuxbus_a vddio vccd0 vssio vccd0 sky130_ef_io__vddio_hvc_clamped_pad
Xgpio0_7_connects gpio0_7_tie_lo_esd gpio0_7_in gpio0_7_tie_hi_esd gpio0_7_enable_vddio
+ gpio0_7_slow gpio0_7_pad_a_esd_0_h gpio0_7_pad_a_esd_1_h gpio0_7_dm[1] gpio0_7_pad_a_noesd_h
+ gpio0_7_analog_en gpio0_7_dm[0] gpio0_7_analog_pol gpio0_7_inp_dis gpio0_7_enable_inp_h
+ gpio0_7_enable_h gpio0_7_hld_h_n gpio0_7_analog_sel gpio0_7_dm[2] gpio0_7_hld_ovr
+ gpio0_7_out gpio0_7_enable_vswitch_h gpio0_7_enable_vdda_h gpio0_7_vtrip_sel gpio0_7_ib_mode_sel
+ gpio0_7_oe_n gpio0_7_in_h gpio0_7_one gpio0_7_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio1_0_connects gpio1_0_one gpio1_0_zero gpio1_0_enable_h gpio1_0_tie_hi_esd gpio1_0_vinref
+ gpio1_0_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xgpio2_2_pad gpio2_2_dm[0] gpio2_2_ib_mode_sel gpio2_2_enable_h gpio2_2_enable_inp_h
+ gpio2_2_slow gpio2_2_vtrip_sel gpio2_2_enable_vddio gpio2_2_enable_vdda_h gpio2_2_pad_a_noesd_h
+ gpio2_2_analog_pol gpio2_2_hld_h_n w_694469_804669# gpio2_2_dm[1] w_692355_801352#
+ gpio2_2_dm[2] w_692253_804670# gpio2_2_pad_a_esd_1_h gpio2_2_tie_hi_esd gpio2_2_enable_vswitch_h
+ gpio2_2_tie_lo_esd gpio2_2_oe_n w_694469_801352# vref_e/amuxbus_b gpio2_2_analog_sel
+ vddio vref_e/amuxbus_a gpio2_2_in_h vddio gpio2_2_inp_dis gpio2_2_out gpio2_2_hld_ovr
+ vccd0 gpio2_2 vccd0 gpio2_2_pad_a_esd_0_h gpio2_2_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio2_2_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio4_5_pad gpio4_5_dm[0] gpio4_5_ib_mode_sel gpio4_5_enable_h gpio4_5_enable_inp_h
+ gpio4_5_slow gpio4_5_vtrip_sel gpio4_5_enable_vddio gpio4_5_enable_vdda_h gpio4_5_pad_a_noesd_h
+ gpio4_5_analog_pol gpio4_5_hld_h_n w_125474_1014469# gpio4_5_dm[1] w_128565_1012355#
+ gpio4_5_dm[2] w_125474_1012253# gpio4_5_pad_a_esd_1_h gpio4_5_tie_hi_esd gpio4_5_enable_vswitch_h
+ gpio4_5_tie_lo_esd gpio4_5_oe_n w_128565_1014469# amuxbus_b_n gpio4_5_analog_sel
+ vddio amuxbus_a_n gpio4_5_in_h vddio gpio4_5_inp_dis gpio4_5_out gpio4_5_hld_ovr
+ vccd0 gpio4_5 vccd0 gpio4_5_pad_a_esd_0_h gpio4_5_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio4_5_in vssd0 sky130_ef_io__gpiov2_pad
Xvcap_e vcap_e_cpos vcap_w/cneg vssio vref_w/vddio_q vddio vcap_w/cneg vccd0 vssa1
+ vccd0 vddio vdda1 vssd0 vref_e/amuxbus_b vref_e/amuxbus_a sky130_fd_io__top_vrefcapv2
Xgpio2_3_connects gpio2_3_tie_lo_esd gpio2_3_in gpio2_3_tie_hi_esd gpio2_3_enable_vddio
+ gpio2_3_slow gpio2_3_pad_a_esd_0_h gpio2_3_pad_a_esd_1_h gpio2_3_dm[1] gpio2_3_pad_a_noesd_h
+ gpio2_3_analog_en gpio2_3_dm[0] gpio2_3_analog_pol gpio2_3_inp_dis gpio2_3_enable_inp_h
+ gpio2_3_enable_h gpio2_3_hld_h_n gpio2_3_analog_sel gpio2_3_dm[2] gpio2_3_hld_ovr
+ gpio2_3_out gpio2_3_enable_vswitch_h gpio2_3_enable_vdda_h gpio2_3_vtrip_sel gpio2_3_ib_mode_sel
+ gpio2_3_oe_n gpio2_3_in_h gpio2_3_one gpio2_3_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xvssa2_0_pad vssd0 vssa2 vddio vssa2_0 vddio vssio vccd0 vdda2 vref_w/vddio_q vref_w/amuxbus_a
+ vref_w/amuxbus_b vcap_w/cneg vccd0 sky130_ef_io__vssa_hvc_clamped_pad
Xgpio3_6_connects gpio3_6_tie_lo_esd gpio3_6_pad_a_esd_1_h gpio3_6_dm[1] gpio3_6_dm[0]
+ gpio3_6_analog_pol gpio3_6_inp_dis gpio3_6_enable_h gpio3_6_hld_h_n gpio3_6_dm[2]
+ gpio3_6_hld_ovr gpio3_6_out gpio3_6_enable_vswitch_h gpio3_6_enable_vdda_h gpio3_6_vtrip_sel
+ gpio3_6_oe_n gpio3_6_tie_hi_esd gpio3_6_in gpio3_6_enable_vddio gpio3_6_slow gpio3_6_pad_a_esd_0_h
+ gpio3_6_pad_a_noesd_h gpio3_6_analog_en gpio3_6_analog_sel gpio3_6_ib_mode_sel gpio3_6_in_h
+ gpio3_6_zero gpio3_6_one gpio3_6_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xvdda2_1_pad vref_w/vddio_q vcap_w/cneg vssio vdda2_1 vref_w/amuxbus_b vref_w/amuxbus_a
+ vdda2 vssd0 vccd0 vssa2 vddio vddio vccd0 sky130_ef_io__vdda_hvc_clamped_pad
Xgpio1_2_pad vcap_w/cneg vddio vssio vssd0 vssa1 vref_w/vddio_q vddio vdda1 vccd0
+ vccd0 gpio1_2 vref_e/amuxbus_a vref_e/amuxbus_b gpio1_2_dm[0] gpio1_2_dm[1] gpio1_2_dm[2]
+ gpio1_2_inp_dis gpio1_2_vtrip_sel gpio1_2_ib_mode_sel[0] gpio1_2_ib_mode_sel[1]
+ gpio1_2_slew_ctl[0] gpio1_2_slew_ctl[1] gpio1_2_hys_trim gpio1_2_hld_ovr gpio1_2_enable_h
+ gpio1_2_hld_h_n gpio1_2_enable_vdda_h gpio1_2_analog_en gpio1_2_enable_inp_h gpio1_2_in
+ gpio1_2_in_h gpio1_0_vinref gpio1_2_out gpio1_2_analog_pol gpio1_2_analog_sel gpio1_2_slow
+ gpio1_2_oe_n gpio1_2_tie_hi_esd gpio1_2_tie_lo_esd gpio1_2_pad_a_esd_0_h gpio1_2_pad_a_esd_1_h
+ gpio1_2_pad_a_noesd_h gpio1_2_enable_vswitch_h gpio1_2_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xgpio5_2_connects gpio5_2_tie_lo_esd gpio5_2_in gpio5_2_tie_hi_esd gpio5_2_enable_vddio
+ gpio5_2_slow gpio5_2_pad_a_esd_0_h gpio5_2_pad_a_esd_1_h gpio5_2_dm[1] gpio5_2_pad_a_noesd_h
+ gpio5_2_analog_en gpio5_2_dm[0] gpio5_2_analog_pol gpio5_2_inp_dis gpio5_2_enable_inp_h
+ gpio5_2_enable_h gpio5_2_hld_h_n gpio5_2_analog_sel gpio5_2_dm[2] gpio5_2_hld_ovr
+ gpio5_2_out gpio5_2_enable_vswitch_h gpio5_2_enable_vdda_h gpio5_2_vtrip_sel gpio5_2_ib_mode_sel
+ gpio5_2_oe_n gpio5_2_in_h gpio5_2_one gpio5_2_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio3_5_pad gpio3_5_dm[0] gpio3_5_ib_mode_sel gpio3_5_enable_h gpio3_5_enable_inp_h
+ gpio3_5_slow gpio3_5_vtrip_sel gpio3_5_enable_vddio gpio3_5_enable_vdda_h gpio3_5_pad_a_noesd_h
+ gpio3_5_analog_pol gpio3_5_hld_h_n w_478474_1014469# gpio3_5_dm[1] w_481565_1012355#
+ gpio3_5_dm[2] w_478474_1012253# gpio3_5_pad_a_esd_1_h gpio3_5_tie_hi_esd gpio3_5_enable_vswitch_h
+ gpio3_5_tie_lo_esd gpio3_5_oe_n w_481565_1014469# amuxbus_b_n gpio3_5_analog_sel
+ vddio amuxbus_a_n gpio3_5_in_h vddio gpio3_5_inp_dis gpio3_5_out gpio3_5_hld_ovr
+ vccd0 gpio3_5 vccd0 gpio3_5_pad_a_esd_0_h gpio3_5_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio3_5_in vssd0 sky130_ef_io__gpiov2_pad
Xvssio_4_pad vdda0 vssd0 vssa0 amuxbus_a_n amuxbus_b_n vssio_4 vref_w/vddio_q vddio
+ vssio vddio vcap_w/cneg vccd0 vccd0 sky130_ef_io__vssio_hvc_clamped_pad
Xgpio6_5_connects gpio6_5_one gpio6_5_zero gpio6_5_enable_h gpio6_5_tie_hi_esd gpio6_7_vinref
+ gpio6_5_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xvssa1_0_pad vssd0 vssa1 vddio vssa1_0 vddio vssio vccd0 vdda1 vref_w/vddio_q vref_e/amuxbus_a
+ vref_e/amuxbus_b vcap_w/cneg vccd0 sky130_ef_io__vssa_hvc_clamped_pad
Xvddio_5_pad vdda2 vcap_w/cneg vddio vref_w/vddio_q vssd0 vddio_5 vssa2 vref_w/amuxbus_b
+ vref_w/amuxbus_a vddio vccd0 vssio vccd0 sky130_ef_io__vddio_hvc_clamped_pad
Xgpio8_1_connects gpio8_1_tie_lo_esd gpio8_1_pad_a_esd_1_h gpio8_1_dm[1] gpio8_1_dm[0]
+ gpio8_1_analog_pol gpio8_1_inp_dis gpio8_1_enable_h gpio8_1_hld_h_n gpio8_1_dm[2]
+ gpio8_1_hld_ovr gpio8_1_out gpio8_1_enable_vswitch_h gpio8_1_enable_vdda_h gpio8_1_vtrip_sel
+ gpio8_1_oe_n gpio8_1_tie_hi_esd gpio8_1_in gpio8_1_enable_vddio gpio8_1_slow gpio8_1_pad_a_esd_0_h
+ gpio8_1_pad_a_noesd_h gpio8_1_analog_en gpio8_1_analog_sel gpio8_1_ib_mode_sel gpio8_1_in_h
+ gpio8_1_zero gpio8_1_one gpio8_1_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xvdda1_1_pad vref_w/vddio_q vcap_w/cneg vssio vdda1_1 vref_e/amuxbus_b vref_e/amuxbus_a
+ vdda1 vssd0 vccd0 vssa1 vddio vddio vccd0 sky130_ef_io__vdda_hvc_clamped_pad
Xgpio0_2_pad gpio0_2_dm[0] gpio0_2_ib_mode_sel gpio0_2_enable_h gpio0_2_enable_inp_h
+ gpio0_2_slow gpio0_2_vtrip_sel gpio0_2_enable_vddio gpio0_2_enable_vdda_h gpio0_2_pad_a_noesd_h
+ gpio0_2_analog_pol gpio0_2_hld_h_n w_694469_120069# gpio0_2_dm[1] w_692355_116752#
+ gpio0_2_dm[2] w_692253_120070# gpio0_2_pad_a_esd_1_h gpio0_2_tie_hi_esd gpio0_2_enable_vswitch_h
+ gpio0_2_tie_lo_esd gpio0_2_oe_n w_694469_116752# vref_e/amuxbus_b gpio0_2_analog_sel
+ vddio vref_e/amuxbus_a gpio0_2_in_h vddio gpio0_2_inp_dis gpio0_2_out gpio0_2_hld_ovr
+ vccd0 gpio0_2 vccd0 gpio0_2_pad_a_esd_0_h gpio0_2_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio0_2_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio2_5_pad gpio2_5_dm[0] gpio2_5_ib_mode_sel gpio2_5_enable_h gpio2_5_enable_inp_h
+ gpio2_5_slow gpio2_5_vtrip_sel gpio2_5_enable_vddio gpio2_5_enable_vdda_h gpio2_5_pad_a_noesd_h
+ gpio2_5_analog_pol gpio2_5_hld_h_n w_694469_887669# gpio2_5_dm[1] w_692355_884352#
+ gpio2_5_dm[2] w_692253_887670# gpio2_5_pad_a_esd_1_h gpio2_5_tie_hi_esd gpio2_5_enable_vswitch_h
+ gpio2_5_tie_lo_esd gpio2_5_oe_n w_694469_884352# vref_e/amuxbus_b gpio2_5_analog_sel
+ vddio vref_e/amuxbus_a gpio2_5_in_h vddio gpio2_5_inp_dis gpio2_5_out gpio2_5_hld_ovr
+ vccd0 gpio2_5 vccd0 gpio2_5_pad_a_esd_0_h gpio2_5_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio2_5_in vssd0 sky130_ef_io__gpiov2_pad
Xvssa0_0_pad vssd0 vssa0 vddio vssa0_0 vddio vssio vccd0 vdda0 vref_w/vddio_q amuxbus_a_n
+ amuxbus_b_n vcap_w/cneg vccd0 sky130_ef_io__vssa_hvc_clamped_pad
Xgpio0_0_connects gpio0_0_tie_lo_esd gpio0_0_in gpio0_0_tie_hi_esd gpio0_0_enable_vddio
+ gpio0_0_slow gpio0_0_pad_a_esd_0_h gpio0_0_pad_a_esd_1_h gpio0_0_dm[1] gpio0_0_pad_a_noesd_h
+ gpio0_0_analog_en gpio0_0_dm[0] gpio0_0_analog_pol gpio0_0_inp_dis gpio0_0_enable_inp_h
+ gpio0_0_enable_h gpio0_0_hld_h_n gpio0_0_analog_sel gpio0_0_dm[2] gpio0_0_hld_ovr
+ gpio0_0_out gpio0_0_enable_vswitch_h gpio0_0_enable_vdda_h gpio0_0_vtrip_sel gpio0_0_ib_mode_sel
+ gpio0_0_oe_n gpio0_0_in_h gpio0_0_one gpio0_0_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio8_1_pad gpio8_1_dm[0] gpio8_1_ib_mode_sel gpio8_1_enable_h gpio8_1_enable_inp_h
+ gpio8_1_slow gpio8_1_vtrip_sel gpio8_1_enable_vddio gpio8_1_enable_vdda_h gpio8_1_pad_a_noesd_h
+ gpio8_1_analog_pol gpio8_1_hld_h_n w_140469_21253# gpio8_1_dm[1] w_137152_23367#
+ gpio8_1_dm[2] w_140469_23367# gpio8_1_pad_a_esd_1_h gpio8_1_tie_hi_esd gpio8_1_enable_vswitch_h
+ gpio8_1_tie_lo_esd gpio8_1_oe_n w_137152_21253# sio_amuxbus_b gpio8_1_analog_sel
+ vddio sio_amuxbus_a gpio8_1_in_h vddio gpio8_1_inp_dis gpio8_1_out gpio8_1_hld_ovr
+ vccd0 gpio8_1 vccd0 gpio8_1_pad_a_esd_0_h gpio8_1_analog_en vssio vdda3 vref_w/vddio_q
+ vcap_w/cneg vssa3 gpio8_1_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio1_3_connects gpio1_3_one gpio1_3_zero gpio1_3_enable_h gpio1_3_tie_hi_esd gpio1_0_vinref
+ gpio1_3_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xgpio2_6_connects gpio2_6_tie_lo_esd gpio2_6_in gpio2_6_tie_hi_esd gpio2_6_enable_vddio
+ gpio2_6_slow gpio2_6_pad_a_esd_0_h gpio2_6_pad_a_esd_1_h gpio2_6_dm[1] gpio2_6_pad_a_noesd_h
+ gpio2_6_analog_en gpio2_6_dm[0] gpio2_6_analog_pol gpio2_6_inp_dis gpio2_6_enable_inp_h
+ gpio2_6_enable_h gpio2_6_hld_h_n gpio2_6_analog_sel gpio2_6_dm[2] gpio2_6_hld_ovr
+ gpio2_6_out gpio2_6_enable_vswitch_h gpio2_6_enable_vdda_h gpio2_6_vtrip_sel gpio2_6_ib_mode_sel
+ gpio2_6_oe_n gpio2_6_in_h gpio2_6_one gpio2_6_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio1_5_pad vcap_w/cneg vddio vssio vssd0 vssa1 vref_w/vddio_q vddio vdda1 vccd0
+ vccd0 gpio1_5 vref_e/amuxbus_a vref_e/amuxbus_b gpio1_5_dm[0] gpio1_5_dm[1] gpio1_5_dm[2]
+ gpio1_5_inp_dis gpio1_5_vtrip_sel gpio1_5_ib_mode_sel[0] gpio1_5_ib_mode_sel[1]
+ gpio1_5_slew_ctl[0] gpio1_5_slew_ctl[1] gpio1_5_hys_trim gpio1_5_hld_ovr gpio1_5_enable_h
+ gpio1_5_hld_h_n gpio1_5_enable_vdda_h gpio1_5_analog_en gpio1_5_enable_inp_h gpio1_5_in
+ gpio1_5_in_h vcap_e_cpos gpio1_5_out gpio1_5_analog_pol gpio1_5_analog_sel gpio1_5_slow
+ gpio1_5_oe_n gpio1_5_tie_hi_esd gpio1_5_tie_lo_esd gpio1_5_pad_a_esd_0_h gpio1_5_pad_a_esd_1_h
+ gpio1_5_pad_a_noesd_h gpio1_5_enable_vswitch_h gpio1_5_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xvssio_7_pad vdda2 vssd0 vssa2 vref_w/amuxbus_a vref_w/amuxbus_b vssio_7 vref_w/vddio_q
+ vddio vssio vddio vcap_w/cneg vccd0 vccd0 sky130_ef_io__vssio_hvc_clamped_pad
Xvccd2_1_pad vdda2 vccd0 vssd2[3] vddio vref_w/amuxbus_b vddio vssio vref_w/amuxbus_a
+ vccd0 vccd2_1 vccd2[3] vssd0 vssa2 vref_w/vddio_q vcap_w/cneg sky130_ef_io__vccd_lvc_clamped3_pad
Xgpio4_2_connects gpio4_2_tie_lo_esd gpio4_2_pad_a_esd_1_h gpio4_2_dm[1] gpio4_2_dm[0]
+ gpio4_2_analog_pol gpio4_2_inp_dis gpio4_2_enable_h gpio4_2_hld_h_n gpio4_2_dm[2]
+ gpio4_2_hld_ovr gpio4_2_out gpio4_2_enable_vswitch_h gpio4_2_enable_vdda_h gpio4_2_vtrip_sel
+ gpio4_2_oe_n gpio4_2_tie_hi_esd gpio4_2_in gpio4_2_enable_vddio gpio4_2_slow gpio4_2_pad_a_esd_0_h
+ gpio4_2_pad_a_noesd_h gpio4_2_analog_en gpio4_2_analog_sel gpio4_2_ib_mode_sel gpio4_2_in_h
+ gpio4_2_zero gpio4_2_one gpio4_2_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio7_1_pad gpio7_1_dm[0] gpio7_1_ib_mode_sel gpio7_1_enable_h gpio7_1_enable_inp_h
+ gpio7_1_slow gpio7_1_vtrip_sel gpio7_1_enable_vddio gpio7_1_enable_vdda_h gpio7_1_pad_a_noesd_h
+ gpio7_1_analog_pol gpio7_1_hld_h_n w_21151_254074# gpio7_1_dm[1] w_23367_257165#
+ gpio7_1_dm[2] w_23367_254074# gpio7_1_pad_a_esd_1_h gpio7_1_tie_hi_esd gpio7_1_enable_vswitch_h
+ gpio7_1_tie_lo_esd gpio7_1_oe_n w_21253_257165# vref_w/amuxbus_b gpio7_1_analog_sel
+ vddio vref_w/amuxbus_a gpio7_1_in_h vddio gpio7_1_inp_dis gpio7_1_out gpio7_1_hld_ovr
+ vccd0 gpio7_1 vccd0 gpio7_1_pad_a_esd_0_h gpio7_1_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio7_1_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio5_5_connects gpio5_5_tie_lo_esd gpio5_5_in gpio5_5_tie_hi_esd gpio5_5_enable_vddio
+ gpio5_5_slow gpio5_5_pad_a_esd_0_h gpio5_5_pad_a_esd_1_h gpio5_5_dm[1] gpio5_5_pad_a_noesd_h
+ gpio5_5_analog_en gpio5_5_dm[0] gpio5_5_analog_pol gpio5_5_inp_dis gpio5_5_enable_inp_h
+ gpio5_5_enable_h gpio5_5_hld_h_n gpio5_5_analog_sel gpio5_5_dm[2] gpio5_5_hld_ovr
+ gpio5_5_out gpio5_5_enable_vswitch_h gpio5_5_enable_vdda_h gpio5_5_vtrip_sel gpio5_5_ib_mode_sel
+ gpio5_5_oe_n gpio5_5_in_h gpio5_5_one gpio5_5_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xvddio_8_pad vdda2 vcap_w/cneg vddio vref_w/vddio_q vssd0 vddio_8 vssa2 vref_w/amuxbus_b
+ vref_w/amuxbus_a vddio vccd0 vssio vccd0 sky130_ef_io__vddio_hvc_clamped_pad
Xresetb_pad resetb_pad_a_esd_h resetb_xres_h_n resetb_filt_in_h resetb_enable_vddio
+ resetb_tie_weak_hi_h resetb_enable_h resetb_pullup_h resetb_en_vddio_sig_h resetb_tie_lo_esd
+ resetb_tie_hi_esd resetb_disable_pullup_h resetb_inp_sel_h vssa3 vssd0 sio_amuxbus_b
+ sio_amuxbus_a vdda3 vccd0 vccd0 vcap_w/cneg vddio vddio vssio resetb vref_w/vddio_q
+ sky130_fd_io__top_xres4v2
Xgpio0_5_pad gpio0_5_dm[0] gpio0_5_ib_mode_sel gpio0_5_enable_h gpio0_5_enable_inp_h
+ gpio0_5_slow gpio0_5_vtrip_sel gpio0_5_enable_vddio gpio0_5_enable_vdda_h gpio0_5_pad_a_noesd_h
+ gpio0_5_analog_pol gpio0_5_hld_h_n w_694469_223069# gpio0_5_dm[1] w_692355_219752#
+ gpio0_5_dm[2] w_692253_223070# gpio0_5_pad_a_esd_1_h gpio0_5_tie_hi_esd gpio0_5_enable_vswitch_h
+ gpio0_5_tie_lo_esd gpio0_5_oe_n w_694469_219752# vref_e/amuxbus_b gpio0_5_analog_sel
+ vddio vref_e/amuxbus_a gpio0_5_in_h vddio gpio0_5_inp_dis gpio0_5_out gpio0_5_hld_ovr
+ vccd0 gpio0_5 vccd0 gpio0_5_pad_a_esd_0_h gpio0_5_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio0_5_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio7_1_connects gpio7_1_tie_lo_esd gpio7_1_in gpio7_1_tie_hi_esd gpio7_1_enable_vddio
+ gpio7_1_slow gpio7_1_pad_a_esd_0_h gpio7_1_pad_a_esd_1_h gpio7_1_dm[1] gpio7_1_pad_a_noesd_h
+ gpio7_1_analog_en gpio7_1_dm[0] gpio7_1_analog_pol gpio7_1_inp_dis gpio7_1_enable_inp_h
+ gpio7_1_enable_h gpio7_1_hld_h_n gpio7_1_analog_sel gpio7_1_dm[2] gpio7_1_hld_ovr
+ gpio7_1_out gpio7_1_enable_vswitch_h gpio7_1_enable_vdda_h gpio7_1_vtrip_sel gpio7_1_ib_mode_sel
+ gpio7_1_oe_n gpio7_1_in_h gpio7_1_one gpio7_1_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xvccd1_1_pad vdda1 vccd0 vssd1[3] vddio vref_e/amuxbus_b vddio vssio vref_e/amuxbus_a
+ vccd0 vccd1_1 vccd1[3] vssd0 vssa1 vref_w/vddio_q vcap_w/cneg sky130_ef_io__vccd_lvc_clamped3_pad
Xgpio6_1_pad vcap_w/cneg vddio vssio vssd0 vssa2 vref_w/vddio_q vddio vdda2 vccd0
+ vccd0 gpio6_1 vref_w/amuxbus_a vref_w/amuxbus_b gpio6_1_dm[0] gpio6_1_dm[1] gpio6_1_dm[2]
+ gpio6_1_inp_dis gpio6_1_vtrip_sel gpio6_1_ib_mode_sel[0] gpio6_1_ib_mode_sel[1]
+ gpio6_1_slew_ctl[0] gpio6_1_slew_ctl[1] gpio6_1_hys_trim gpio6_1_hld_ovr gpio6_1_enable_h
+ gpio6_1_hld_h_n gpio6_1_enable_vdda_h gpio6_1_analog_en gpio6_1_enable_inp_h gpio6_1_in
+ gpio6_1_in_h vcap_w_cpos gpio6_1_out gpio6_1_analog_pol gpio6_1_analog_sel gpio6_1_slow
+ gpio6_1_oe_n gpio6_1_tie_hi_esd gpio6_1_tie_lo_esd gpio6_1_pad_a_esd_0_h gpio6_1_pad_a_esd_1_h
+ gpio6_1_pad_a_noesd_h gpio6_1_enable_vswitch_h gpio6_1_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xgpio8_4_connects gpio8_4_tie_lo_esd gpio8_4_pad_a_esd_1_h gpio8_4_dm[1] gpio8_4_dm[0]
+ gpio8_4_analog_pol gpio8_4_inp_dis gpio8_4_enable_h gpio8_4_hld_h_n gpio8_4_dm[2]
+ gpio8_4_hld_ovr gpio8_4_out gpio8_4_enable_vswitch_h gpio8_4_enable_vdda_h gpio8_4_vtrip_sel
+ gpio8_4_oe_n gpio8_4_tie_hi_esd gpio8_4_in gpio8_4_enable_vddio gpio8_4_slow gpio8_4_pad_a_esd_0_h
+ gpio8_4_pad_a_noesd_h gpio8_4_analog_en gpio8_4_analog_sel gpio8_4_ib_mode_sel gpio8_4_in_h
+ gpio8_4_zero gpio8_4_one gpio8_4_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio8_4_pad gpio8_4_dm[0] gpio8_4_ib_mode_sel gpio8_4_enable_h gpio8_4_enable_inp_h
+ gpio8_4_slow gpio8_4_vtrip_sel gpio8_4_enable_vddio gpio8_4_enable_vdda_h gpio8_4_pad_a_noesd_h
+ gpio8_4_analog_pol gpio8_4_hld_h_n w_389469_21253# gpio8_4_dm[1] w_386152_23367#
+ gpio8_4_dm[2] w_389469_23367# gpio8_4_pad_a_esd_1_h gpio8_4_tie_hi_esd gpio8_4_enable_vswitch_h
+ gpio8_4_tie_lo_esd gpio8_4_oe_n w_386152_21253# sio_amuxbus_b gpio8_4_analog_sel
+ vddio sio_amuxbus_a gpio8_4_in_h vddio gpio8_4_inp_dis gpio8_4_out gpio8_4_hld_ovr
+ vccd0 gpio8_4 vccd0 gpio8_4_pad_a_esd_0_h gpio8_4_analog_en vssio vdda3 vref_w/vddio_q
+ vcap_w/cneg vssa3 gpio8_4_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio0_3_connects gpio0_3_tie_lo_esd gpio0_3_in gpio0_3_tie_hi_esd gpio0_3_enable_vddio
+ gpio0_3_slow gpio0_3_pad_a_esd_0_h gpio0_3_pad_a_esd_1_h gpio0_3_dm[1] gpio0_3_pad_a_noesd_h
+ gpio0_3_analog_en gpio0_3_dm[0] gpio0_3_analog_pol gpio0_3_inp_dis gpio0_3_enable_inp_h
+ gpio0_3_enable_h gpio0_3_hld_h_n gpio0_3_analog_sel gpio0_3_dm[2] gpio0_3_hld_ovr
+ gpio0_3_out gpio0_3_enable_vswitch_h gpio0_3_enable_vdda_h gpio0_3_vtrip_sel gpio0_3_ib_mode_sel
+ gpio0_3_oe_n gpio0_3_in_h gpio0_3_one gpio0_3_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xvccd0_1_pad vdda3 vccd0 sio_amuxbus_b sio_amuxbus_a vccd0_1 vccd0 vddio vssd0 vssio
+ vssa3 vddio vref_w/vddio_q vcap_w/cneg sky130_ef_io__vccd_lvc_clamped_pad
Xgpio5_1_pad gpio5_1_dm[0] gpio5_1_ib_mode_sel gpio5_1_enable_h gpio5_1_enable_inp_h
+ gpio5_1_slow gpio5_1_vtrip_sel gpio5_1_enable_vddio gpio5_1_enable_vdda_h gpio5_1_pad_a_noesd_h
+ gpio5_1_analog_pol gpio5_1_hld_h_n w_21151_916674# gpio5_1_dm[1] w_23367_919765#
+ gpio5_1_dm[2] w_23367_916674# gpio5_1_pad_a_esd_1_h gpio5_1_tie_hi_esd gpio5_1_enable_vswitch_h
+ gpio5_1_tie_lo_esd gpio5_1_oe_n w_21253_919765# vref_w/amuxbus_b gpio5_1_analog_sel
+ vddio vref_w/amuxbus_a gpio5_1_in_h vddio gpio5_1_inp_dis gpio5_1_out gpio5_1_hld_ovr
+ vccd0 gpio5_1 vccd0 gpio5_1_pad_a_esd_0_h gpio5_1_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio5_1_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio1_6_connects gpio1_6_one gpio1_6_zero gpio1_6_enable_h gpio1_6_tie_hi_esd vcap_e_cpos
+ gpio1_6_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xgpio7_4_pad gpio7_4_dm[0] gpio7_4_ib_mode_sel gpio7_4_enable_h gpio7_4_enable_inp_h
+ gpio7_4_slow gpio7_4_vtrip_sel gpio7_4_enable_vddio gpio7_4_enable_vdda_h gpio7_4_pad_a_noesd_h
+ gpio7_4_analog_pol gpio7_4_hld_h_n w_21151_148074# gpio7_4_dm[1] w_23367_151165#
+ gpio7_4_dm[2] w_23367_148074# gpio7_4_pad_a_esd_1_h gpio7_4_tie_hi_esd gpio7_4_enable_vswitch_h
+ gpio7_4_tie_lo_esd gpio7_4_oe_n w_21253_151165# vref_w/amuxbus_b gpio7_4_analog_sel
+ vddio vref_w/amuxbus_a gpio7_4_in_h vddio gpio7_4_inp_dis gpio7_4_out gpio7_4_hld_ovr
+ vccd0 gpio7_4 vccd0 gpio7_4_pad_a_esd_0_h gpio7_4_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio7_4_in vssd0 sky130_ef_io__gpiov2_pad
Xvref_e vref_e_ref_sel[4] vref_e_ref_sel[3] vref_e_ref_sel[1] vref_e_vrefgen_en vref_e_hld_h_n
+ vref_e_enable_h vref_e_ref_sel[2] vref_e_ref_sel[0] gpio1_0_vinref vref_w/vddio_q
+ vddio vssio vssa1 vccd0 vccd0 vddio vcap_w/cneg vdda1 vssd0 vref_e/amuxbus_b vref_e/amuxbus_a
+ sky130_fd_io__top_gpiovrefv2
Xgpio3_2_connects gpio3_2_tie_lo_esd gpio3_2_pad_a_esd_1_h gpio3_2_dm[1] gpio3_2_dm[0]
+ gpio3_2_analog_pol gpio3_2_inp_dis gpio3_2_enable_h gpio3_2_hld_h_n gpio3_2_dm[2]
+ gpio3_2_hld_ovr gpio3_2_out gpio3_2_enable_vswitch_h gpio3_2_enable_vdda_h gpio3_2_vtrip_sel
+ gpio3_2_oe_n gpio3_2_tie_hi_esd gpio3_2_in gpio3_2_enable_vddio gpio3_2_slow gpio3_2_pad_a_esd_0_h
+ gpio3_2_pad_a_noesd_h gpio3_2_analog_en gpio3_2_analog_sel gpio3_2_ib_mode_sel gpio3_2_in_h
+ gpio3_2_zero gpio3_2_one gpio3_2_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio4_5_connects gpio4_5_tie_lo_esd gpio4_5_pad_a_esd_1_h gpio4_5_dm[1] gpio4_5_dm[0]
+ gpio4_5_analog_pol gpio4_5_inp_dis gpio4_5_enable_h gpio4_5_hld_h_n gpio4_5_dm[2]
+ gpio4_5_hld_ovr gpio4_5_out gpio4_5_enable_vswitch_h gpio4_5_enable_vdda_h gpio4_5_vtrip_sel
+ gpio4_5_oe_n gpio4_5_tie_hi_esd gpio4_5_in gpio4_5_enable_vddio gpio4_5_slow gpio4_5_pad_a_esd_0_h
+ gpio4_5_pad_a_noesd_h gpio4_5_analog_en gpio4_5_analog_sel gpio4_5_ib_mode_sel gpio4_5_in_h
+ gpio4_5_zero gpio4_5_one gpio4_5_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio4_1_pad gpio4_1_dm[0] gpio4_1_ib_mode_sel gpio4_1_enable_h gpio4_1_enable_inp_h
+ gpio4_1_slow gpio4_1_vtrip_sel gpio4_1_enable_vddio gpio4_1_enable_vdda_h gpio4_1_pad_a_noesd_h
+ gpio4_1_analog_pol gpio4_1_hld_h_n w_267474_1014469# gpio4_1_dm[1] w_270565_1012355#
+ gpio4_1_dm[2] w_267474_1012253# gpio4_1_pad_a_esd_1_h gpio4_1_tie_hi_esd gpio4_1_enable_vswitch_h
+ gpio4_1_tie_lo_esd gpio4_1_oe_n w_270565_1014469# amuxbus_b_n gpio4_1_analog_sel
+ vddio amuxbus_a_n gpio4_1_in_h vddio gpio4_1_inp_dis gpio4_1_out gpio4_1_hld_ovr
+ vccd0 gpio4_1 vccd0 gpio4_1_pad_a_esd_0_h gpio4_1_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio4_1_in vssd0 sky130_ef_io__gpiov2_pad
Xmuxsplit_sw vref_w/amuxbus_a sio_amuxbus_a vref_w/amuxbus_b sio_amuxbus_b muxsplit_sw_enable_vdda_h
+ muxsplit_sw_hld_vdda_h_n muxsplit_sw_switch_aa_s0 muxsplit_sw_switch_aa_sl muxsplit_sw_switch_aa_sr
+ muxsplit_sw_switch_bb_s0 muxsplit_sw_switch_bb_sl muxsplit_sw_switch_bb_sr vssd0
+ vssio vddio vccd0 vref_w/vddio_q vddio vccd0 w_4981_42974# w_11281_42974# vdda3
+ vssa3 vcap_w/cneg sky130_fd_io__top_amuxsplitv2
Xvssd2_1_pad vdda2 vcap_w/cneg vssd2[2] vccd0 vssd0 vssa2 vref_w/amuxbus_b vref_w/amuxbus_a
+ vssd2_1 vddio vddio vccd0 vref_w/vddio_q vssio vccd2[2] sky130_ef_io__vssd_lvc_clamped3_pad
Xgpio6_4_pad vcap_w/cneg vddio vssio vssd0 vssa2 vref_w/vddio_q vddio vdda2 vccd0
+ vccd0 gpio6_4 vref_w/amuxbus_a vref_w/amuxbus_b gpio6_4_dm[0] gpio6_4_dm[1] gpio6_4_dm[2]
+ gpio6_4_inp_dis gpio6_4_vtrip_sel gpio6_4_ib_mode_sel[0] gpio6_4_ib_mode_sel[1]
+ gpio6_4_slew_ctl[0] gpio6_4_slew_ctl[1] gpio6_4_hys_trim gpio6_4_hld_ovr gpio6_4_enable_h
+ gpio6_4_hld_h_n gpio6_4_enable_vdda_h gpio6_4_analog_en gpio6_4_enable_inp_h gpio6_4_in
+ gpio6_4_in_h gpio6_7_vinref gpio6_4_out gpio6_4_analog_pol gpio6_4_analog_sel gpio6_4_slow
+ gpio6_4_oe_n gpio6_4_tie_hi_esd gpio6_4_tie_lo_esd gpio6_4_pad_a_esd_0_h gpio6_4_pad_a_esd_1_h
+ gpio6_4_pad_a_noesd_h gpio6_4_enable_vswitch_h gpio6_4_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xgpio6_1_connects gpio6_1_one gpio6_1_zero gpio6_1_enable_h gpio6_1_tie_hi_esd vcap_w_cpos
+ gpio6_1_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xgpio8_7_pad gpio8_7_dm[0] gpio8_7_ib_mode_sel gpio8_7_enable_h gpio8_7_enable_inp_h
+ gpio8_7_slow gpio8_7_vtrip_sel gpio8_7_enable_vddio gpio8_7_enable_vdda_h gpio8_7_pad_a_noesd_h
+ gpio8_7_analog_pol gpio8_7_hld_h_n w_458469_21253# gpio8_7_dm[1] w_455152_23367#
+ gpio8_7_dm[2] w_458469_23367# gpio8_7_pad_a_esd_1_h gpio8_7_tie_hi_esd gpio8_7_enable_vswitch_h
+ gpio8_7_tie_lo_esd gpio8_7_oe_n w_455152_21253# sio_amuxbus_b gpio8_7_analog_sel
+ vddio sio_amuxbus_a gpio8_7_in_h vddio gpio8_7_inp_dis gpio8_7_out gpio8_7_hld_ovr
+ vccd0 gpio8_7 vccd0 gpio8_7_pad_a_esd_0_h gpio8_7_analog_en vssio vdda3 vref_w/vddio_q
+ vcap_w/cneg vssa3 gpio8_7_in vssd0 sky130_ef_io__gpiov2_pad
Xpwrdet_s pwrdet_in1_vddd_hv pwrdet_in2_vddd_hv pwrdet_out3_vddio_hv pwrdet_out1_vddio_hv
+ pwrdet_out2_vddio_hv pwrdet_out2_vddd_hv pwrdet_out1_vddd_hv pwrdet_in1_vddio_hv
+ pwrdet_vddio_present_vddd_hv pwrdet_vddd_present_vddio_hv pwrdet_tie_lo_esd pwrdet_rst_por_hv_n
+ pwrdet_out3_vddd_hv pwrdet_in3_vddio_hv pwrdet_in2_vddio_hv pwrdet_in3_vddd_hv pwrdet_s/vssio_q
+ vccd0 vdda3 vssa3 vref_w/vddio_q vdda3 vssd0 sky130_fd_io__top_pwrdetv2
Xgpio7_4_connects gpio7_4_tie_lo_esd gpio7_4_in gpio7_4_tie_hi_esd gpio7_4_enable_vddio
+ gpio7_4_slow gpio7_4_pad_a_esd_0_h gpio7_4_pad_a_esd_1_h gpio7_4_dm[1] gpio7_4_pad_a_noesd_h
+ gpio7_4_analog_en gpio7_4_dm[0] gpio7_4_analog_pol gpio7_4_inp_dis gpio7_4_enable_inp_h
+ gpio7_4_enable_h gpio7_4_hld_h_n gpio7_4_analog_sel gpio7_4_dm[2] gpio7_4_hld_ovr
+ gpio7_4_out gpio7_4_enable_vswitch_h gpio7_4_enable_vdda_h gpio7_4_vtrip_sel gpio7_4_ib_mode_sel
+ gpio7_4_oe_n gpio7_4_in_h gpio7_4_one gpio7_4_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio8_7_connects gpio8_7_tie_lo_esd gpio8_7_pad_a_esd_1_h gpio8_7_dm[1] gpio8_7_dm[0]
+ gpio8_7_analog_pol gpio8_7_inp_dis gpio8_7_enable_h gpio8_7_hld_h_n gpio8_7_dm[2]
+ gpio8_7_hld_ovr gpio8_7_out gpio8_7_enable_vswitch_h gpio8_7_enable_vdda_h gpio8_7_vtrip_sel
+ gpio8_7_oe_n gpio8_7_tie_hi_esd gpio8_7_in gpio8_7_enable_vddio gpio8_7_slow gpio8_7_pad_a_esd_0_h
+ gpio8_7_pad_a_noesd_h gpio8_7_analog_en gpio8_7_analog_sel gpio8_7_ib_mode_sel gpio8_7_in_h
+ gpio8_7_zero gpio8_7_one gpio8_7_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio3_1_pad gpio3_1_dm[0] gpio3_1_ib_mode_sel gpio3_1_enable_h gpio3_1_enable_inp_h
+ gpio3_1_slow gpio3_1_vtrip_sel gpio3_1_enable_vddio gpio3_1_enable_vdda_h gpio3_1_pad_a_noesd_h
+ gpio3_1_analog_pol gpio3_1_hld_h_n w_620474_1014469# gpio3_1_dm[1] w_623565_1012355#
+ gpio3_1_dm[2] w_620474_1012253# gpio3_1_pad_a_esd_1_h gpio3_1_tie_hi_esd gpio3_1_enable_vswitch_h
+ gpio3_1_tie_lo_esd gpio3_1_oe_n w_623565_1014469# amuxbus_b_n gpio3_1_analog_sel
+ vddio amuxbus_a_n gpio3_1_in_h vddio gpio3_1_inp_dis gpio3_1_out gpio3_1_hld_ovr
+ vccd0 gpio3_1 vccd0 gpio3_1_pad_a_esd_0_h gpio3_1_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio3_1_in vssd0 sky130_ef_io__gpiov2_pad
Xvssio_0_pad vdda1 vssd0 vssa1 vref_e/amuxbus_a vref_e/amuxbus_b vssio_0 vref_w/vddio_q
+ vddio vssio vddio vcap_w/cneg vccd0 vccd0 sky130_ef_io__vssio_hvc_clamped_pad
Xvssd1_1_pad vdda1 vcap_w/cneg vssd1[2] vccd0 vssd0 vssa1 vref_e/amuxbus_b vref_e/amuxbus_a
+ vssd1_1 vddio vddio vccd0 vref_w/vddio_q vssio vccd1[2] sky130_ef_io__vssd_lvc_clamped3_pad
Xgpio5_4_pad gpio5_4_dm[0] gpio5_4_ib_mode_sel gpio5_4_enable_h gpio5_4_enable_inp_h
+ gpio5_4_slow gpio5_4_vtrip_sel gpio5_4_enable_vddio gpio5_4_enable_vdda_h gpio5_4_pad_a_noesd_h
+ gpio5_4_analog_pol gpio5_4_hld_h_n w_21151_833674# gpio5_4_dm[1] w_23367_836765#
+ gpio5_4_dm[2] w_23367_833674# gpio5_4_pad_a_esd_1_h gpio5_4_tie_hi_esd gpio5_4_enable_vswitch_h
+ gpio5_4_tie_lo_esd gpio5_4_oe_n w_21253_836765# vref_w/amuxbus_b gpio5_4_analog_sel
+ vddio vref_w/amuxbus_a gpio5_4_in_h vddio gpio5_4_inp_dis gpio5_4_out gpio5_4_hld_ovr
+ vccd0 gpio5_4 vccd0 gpio5_4_pad_a_esd_0_h gpio5_4_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio5_4_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio7_7_pad gpio7_7_dm[0] gpio7_7_ib_mode_sel gpio7_7_enable_h gpio7_7_enable_inp_h
+ gpio7_7_slow gpio7_7_vtrip_sel gpio7_7_enable_vddio gpio7_7_enable_vdda_h gpio7_7_pad_a_noesd_h
+ gpio7_7_analog_pol gpio7_7_hld_h_n w_21151_85074# gpio7_7_dm[1] w_23367_88165# gpio7_7_dm[2]
+ w_23367_85074# gpio7_7_pad_a_esd_1_h gpio7_7_tie_hi_esd gpio7_7_enable_vswitch_h
+ gpio7_7_tie_lo_esd gpio7_7_oe_n w_21253_88165# vref_w/amuxbus_b gpio7_7_analog_sel
+ vddio vref_w/amuxbus_a gpio7_7_in_h vddio gpio7_7_inp_dis gpio7_7_out gpio7_7_hld_ovr
+ vccd0 gpio7_7 vccd0 gpio7_7_pad_a_esd_0_h gpio7_7_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio7_7_in vssd0 sky130_ef_io__gpiov2_pad
Xvddio_1_pad vdda1 vcap_w/cneg vddio vref_w/vddio_q vssd0 vddio_1 vssa1 vref_e/amuxbus_b
+ vref_e/amuxbus_a vddio vccd0 vssio vccd0 sky130_ef_io__vddio_hvc_clamped_pad
Xgpio0_6_connects gpio0_6_tie_lo_esd gpio0_6_in gpio0_6_tie_hi_esd gpio0_6_enable_vddio
+ gpio0_6_slow gpio0_6_pad_a_esd_0_h gpio0_6_pad_a_esd_1_h gpio0_6_dm[1] gpio0_6_pad_a_noesd_h
+ gpio0_6_analog_en gpio0_6_dm[0] gpio0_6_analog_pol gpio0_6_inp_dis gpio0_6_enable_inp_h
+ gpio0_6_enable_h gpio0_6_hld_h_n gpio0_6_analog_sel gpio0_6_dm[2] gpio0_6_hld_ovr
+ gpio0_6_out gpio0_6_enable_vswitch_h gpio0_6_enable_vdda_h gpio0_6_vtrip_sel gpio0_6_ib_mode_sel
+ gpio0_6_oe_n gpio0_6_in_h gpio0_6_one gpio0_6_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xvdda3_0_pad vref_w/vddio_q vcap_w/cneg vssio vdda3_0 sio_amuxbus_b sio_amuxbus_a
+ vdda3 vssd0 vccd0 vssa3 vddio vddio vccd0 sky130_ef_io__vdda_hvc_clamped_pad
Xgpio2_1_pad gpio2_1_dm[0] gpio2_1_ib_mode_sel gpio2_1_enable_h gpio2_1_enable_inp_h
+ gpio2_1_slow gpio2_1_vtrip_sel gpio2_1_enable_vddio gpio2_1_enable_vdda_h gpio2_1_pad_a_noesd_h
+ gpio2_1_analog_pol gpio2_1_hld_h_n w_694469_783669# gpio2_1_dm[1] w_692355_780352#
+ gpio2_1_dm[2] w_692253_783670# gpio2_1_pad_a_esd_1_h gpio2_1_tie_hi_esd gpio2_1_enable_vswitch_h
+ gpio2_1_tie_lo_esd gpio2_1_oe_n w_694469_780352# vref_e/amuxbus_b gpio2_1_analog_sel
+ vddio vref_e/amuxbus_a gpio2_1_in_h vddio gpio2_1_inp_dis gpio2_1_out gpio2_1_hld_ovr
+ vccd0 gpio2_1 vccd0 gpio2_1_pad_a_esd_0_h gpio2_1_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio2_1_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio2_2_connects gpio2_2_tie_lo_esd gpio2_2_in gpio2_2_tie_hi_esd gpio2_2_enable_vddio
+ gpio2_2_slow gpio2_2_pad_a_esd_0_h gpio2_2_pad_a_esd_1_h gpio2_2_dm[1] gpio2_2_pad_a_noesd_h
+ gpio2_2_analog_en gpio2_2_dm[0] gpio2_2_analog_pol gpio2_2_inp_dis gpio2_2_enable_inp_h
+ gpio2_2_enable_h gpio2_2_hld_h_n gpio2_2_analog_sel gpio2_2_dm[2] gpio2_2_hld_ovr
+ gpio2_2_out gpio2_2_enable_vswitch_h gpio2_2_enable_vdda_h gpio2_2_vtrip_sel gpio2_2_ib_mode_sel
+ gpio2_2_oe_n gpio2_2_in_h gpio2_2_one gpio2_2_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio4_4_pad gpio4_4_dm[0] gpio4_4_ib_mode_sel gpio4_4_enable_h gpio4_4_enable_inp_h
+ gpio4_4_slow gpio4_4_vtrip_sel gpio4_4_enable_vddio gpio4_4_enable_vdda_h gpio4_4_pad_a_noesd_h
+ gpio4_4_analog_pol gpio4_4_hld_h_n w_149474_1014469# gpio4_4_dm[1] w_152565_1012355#
+ gpio4_4_dm[2] w_149474_1012253# gpio4_4_pad_a_esd_1_h gpio4_4_tie_hi_esd gpio4_4_enable_vswitch_h
+ gpio4_4_tie_lo_esd gpio4_4_oe_n w_152565_1014469# amuxbus_b_n gpio4_4_analog_sel
+ vddio amuxbus_a_n gpio4_4_in_h vddio gpio4_4_inp_dis gpio4_4_out gpio4_4_hld_ovr
+ vccd0 gpio4_4 vccd0 gpio4_4_pad_a_esd_0_h gpio4_4_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio4_4_in vssd0 sky130_ef_io__gpiov2_pad
Xvssd0_1_pad vdda3 vssd0_1 vccd0 vddio vddio sio_amuxbus_a sio_amuxbus_b vref_w/vddio_q
+ vssd0 vssio vcap_w/cneg vccd0 vssa3 sky130_ef_io__vssd_lvc_clamped_pad
Xselect_pad select_dm[0] select_ib_mode_sel select_enable_h select_enable_inp_h select_slow
+ select_vtrip_sel select_enable_vddio select_enable_vdda_h select_pad_a_noesd_h select_analog_pol
+ select_hld_h_n w_72469_21253# select_dm[1] w_69152_23367# select_dm[2] w_72469_23367#
+ select_pad_a_esd_1_h select_tie_hi_esd select_enable_vswitch_h select_tie_lo_esd
+ select_oe_n w_69152_21253# sio_amuxbus_b select_analog_sel vddio sio_amuxbus_a select_in_h
+ vddio select_inp_dis select_out select_hld_ovr vccd0 select vccd0 select_pad_a_esd_0_h
+ select_analog_en vssio vdda3 vref_w/vddio_q vcap_w/cneg vssa3 select_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio3_5_connects gpio3_5_tie_lo_esd gpio3_5_pad_a_esd_1_h gpio3_5_dm[1] gpio3_5_dm[0]
+ gpio3_5_analog_pol gpio3_5_inp_dis gpio3_5_enable_h gpio3_5_hld_h_n gpio3_5_dm[2]
+ gpio3_5_hld_ovr gpio3_5_out gpio3_5_enable_vswitch_h gpio3_5_enable_vdda_h gpio3_5_vtrip_sel
+ gpio3_5_oe_n gpio3_5_tie_hi_esd gpio3_5_in gpio3_5_enable_vddio gpio3_5_slow gpio3_5_pad_a_esd_0_h
+ gpio3_5_pad_a_noesd_h gpio3_5_analog_en gpio3_5_analog_sel gpio3_5_ib_mode_sel gpio3_5_in_h
+ gpio3_5_zero gpio3_5_one gpio3_5_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio6_7_pad vcap_w/cneg vddio vssio vssd0 vssa2 vref_w/vddio_q vddio vdda2 vccd0
+ vccd0 gpio6_7 vref_w/amuxbus_a vref_w/amuxbus_b gpio6_7_dm[0] gpio6_7_dm[1] gpio6_7_dm[2]
+ gpio6_7_inp_dis gpio6_7_vtrip_sel gpio6_7_ib_mode_sel[0] gpio6_7_ib_mode_sel[1]
+ gpio6_7_slew_ctl[0] gpio6_7_slew_ctl[1] gpio6_7_hys_trim gpio6_7_hld_ovr gpio6_7_enable_h
+ gpio6_7_hld_h_n gpio6_7_enable_vdda_h gpio6_7_analog_en gpio6_7_enable_inp_h gpio6_7_in
+ gpio6_7_in_h gpio6_7_vinref gpio6_7_out gpio6_7_analog_pol gpio6_7_analog_sel gpio6_7_slow
+ gpio6_7_oe_n gpio6_7_tie_hi_esd gpio6_7_tie_lo_esd gpio6_7_pad_a_esd_0_h gpio6_7_pad_a_esd_1_h
+ gpio6_7_pad_a_noesd_h gpio6_7_enable_vswitch_h gpio6_7_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xxi1_pad vccd0 vref_w/vddio_q vccd0 vcap_w/cneg vssd0 sio_amuxbus_b sio_amuxbus_a
+ xi1_core vssa3 vddio vddio vdda3 vssio xi1 sky130_fd_io__top_analog_pad
Xgpio5_1_connects gpio5_1_tie_lo_esd gpio5_1_in gpio5_1_tie_hi_esd gpio5_1_enable_vddio
+ gpio5_1_slow gpio5_1_pad_a_esd_0_h gpio5_1_pad_a_esd_1_h gpio5_1_dm[1] gpio5_1_pad_a_noesd_h
+ gpio5_1_analog_en gpio5_1_dm[0] gpio5_1_analog_pol gpio5_1_inp_dis gpio5_1_enable_inp_h
+ gpio5_1_enable_h gpio5_1_hld_h_n gpio5_1_analog_sel gpio5_1_dm[2] gpio5_1_hld_ovr
+ gpio5_1_out gpio5_1_enable_vswitch_h gpio5_1_enable_vdda_h gpio5_1_vtrip_sel gpio5_1_ib_mode_sel
+ gpio5_1_oe_n gpio5_1_in_h gpio5_1_one gpio5_1_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio1_1_pad vcap_w/cneg vddio vssio vssd0 vssa1 vref_w/vddio_q vddio vdda1 vccd0
+ vccd0 gpio1_1 vref_e/amuxbus_a vref_e/amuxbus_b gpio1_1_dm[0] gpio1_1_dm[1] gpio1_1_dm[2]
+ gpio1_1_inp_dis gpio1_1_vtrip_sel gpio1_1_ib_mode_sel[0] gpio1_1_ib_mode_sel[1]
+ gpio1_1_slew_ctl[0] gpio1_1_slew_ctl[1] gpio1_1_hys_trim gpio1_1_hld_ovr gpio1_1_enable_h
+ gpio1_1_hld_h_n gpio1_1_enable_vdda_h gpio1_1_analog_en gpio1_1_enable_inp_h gpio1_1_in
+ gpio1_1_in_h gpio1_0_vinref gpio1_1_out gpio1_1_analog_pol gpio1_1_analog_sel gpio1_1_slow
+ gpio1_1_oe_n gpio1_1_tie_hi_esd gpio1_1_tie_lo_esd gpio1_1_pad_a_esd_0_h gpio1_1_pad_a_esd_1_h
+ gpio1_1_pad_a_noesd_h gpio1_1_enable_vswitch_h gpio1_1_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xvdda2_0_pad vref_w/vddio_q vcap_w/cneg vssio vdda2_0 vref_w/amuxbus_b vref_w/amuxbus_a
+ vdda2 vssd0 vccd0 vssa2 vddio vddio vccd0 sky130_ef_io__vdda_hvc_clamped_pad
Xgpio6_4_connects gpio6_4_one gpio6_4_zero gpio6_4_enable_h gpio6_4_tie_hi_esd gpio6_7_vinref
+ gpio6_4_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xvssio_3_pad vdda0 vssd0 vssa0 amuxbus_a_n amuxbus_b_n vssio_3 vref_w/vddio_q vddio
+ vssio vddio vcap_w/cneg vccd0 vccd0 sky130_ef_io__vssio_hvc_clamped_pad
Xgpio3_4_pad gpio3_4_dm[0] gpio3_4_ib_mode_sel gpio3_4_enable_h gpio3_4_enable_inp_h
+ gpio3_4_slow gpio3_4_vtrip_sel gpio3_4_enable_vddio gpio3_4_enable_vdda_h gpio3_4_pad_a_noesd_h
+ gpio3_4_analog_pol gpio3_4_hld_h_n w_502474_1014469# gpio3_4_dm[1] w_505565_1012355#
+ gpio3_4_dm[2] w_502474_1012253# gpio3_4_pad_a_esd_1_h gpio3_4_tie_hi_esd gpio3_4_enable_vswitch_h
+ gpio3_4_tie_lo_esd gpio3_4_oe_n w_505565_1014469# amuxbus_b_n gpio3_4_analog_sel
+ vddio amuxbus_a_n gpio3_4_in_h vddio gpio3_4_inp_dis gpio3_4_out gpio3_4_hld_ovr
+ vccd0 gpio3_4 vccd0 gpio3_4_pad_a_esd_0_h gpio3_4_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio3_4_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio7_7_connects gpio7_7_tie_lo_esd gpio7_7_in gpio7_7_tie_hi_esd gpio7_7_enable_vddio
+ gpio7_7_slow gpio7_7_pad_a_esd_0_h gpio7_7_pad_a_esd_1_h gpio7_7_dm[1] gpio7_7_pad_a_noesd_h
+ gpio7_7_analog_en gpio7_7_dm[0] gpio7_7_analog_pol gpio7_7_inp_dis gpio7_7_enable_inp_h
+ gpio7_7_enable_h gpio7_7_hld_h_n gpio7_7_analog_sel gpio7_7_dm[2] gpio7_7_hld_ovr
+ gpio7_7_out gpio7_7_enable_vswitch_h gpio7_7_enable_vdda_h gpio7_7_vtrip_sel gpio7_7_ib_mode_sel
+ gpio7_7_oe_n gpio7_7_in_h gpio7_7_one gpio7_7_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio5_7_pad gpio5_7_dm[0] gpio5_7_ib_mode_sel gpio5_7_enable_h gpio5_7_enable_inp_h
+ gpio5_7_slow gpio5_7_vtrip_sel gpio5_7_enable_vddio gpio5_7_enable_vdda_h gpio5_7_pad_a_noesd_h
+ gpio5_7_analog_pol gpio5_7_hld_h_n w_21151_770674# gpio5_7_dm[1] w_23367_773765#
+ gpio5_7_dm[2] w_23367_770674# gpio5_7_pad_a_esd_1_h gpio5_7_tie_hi_esd gpio5_7_enable_vswitch_h
+ gpio5_7_tie_lo_esd gpio5_7_oe_n w_21253_773765# vref_w/amuxbus_b gpio5_7_analog_sel
+ vddio vref_w/amuxbus_a gpio5_7_in_h vddio gpio5_7_inp_dis gpio5_7_out gpio5_7_hld_ovr
+ vccd0 gpio5_7 vccd0 gpio5_7_pad_a_esd_0_h gpio5_7_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio5_7_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio8_0_connects gpio8_0_tie_lo_esd gpio8_0_pad_a_esd_1_h gpio8_0_dm[1] gpio8_0_dm[0]
+ gpio8_0_analog_pol gpio8_0_inp_dis gpio8_0_enable_h gpio8_0_hld_h_n gpio8_0_dm[2]
+ gpio8_0_hld_ovr gpio8_0_out gpio8_0_enable_vswitch_h gpio8_0_enable_vdda_h gpio8_0_vtrip_sel
+ gpio8_0_oe_n gpio8_0_tie_hi_esd gpio8_0_in gpio8_0_enable_vddio gpio8_0_slow gpio8_0_pad_a_esd_0_h
+ gpio8_0_pad_a_noesd_h gpio8_0_analog_en gpio8_0_analog_sel gpio8_0_ib_mode_sel gpio8_0_in_h
+ gpio8_0_zero gpio8_0_one gpio8_0_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xvddio_4_pad vdda0 vcap_w/cneg vddio vref_w/vddio_q vssd0 vddio_4 vssa0 amuxbus_b_n
+ amuxbus_a_n vddio vccd0 vssio vccd0 sky130_ef_io__vddio_hvc_clamped_pad
Xmuxsplit_nw amuxbus_a_n vref_w/amuxbus_a amuxbus_b_n vref_w/amuxbus_b muxsplit_nw_enable_vdda_h
+ muxsplit_nw_hld_vdda_h_n muxsplit_nw_switch_aa_s0 muxsplit_nw_switch_aa_sl muxsplit_nw_switch_aa_sr
+ muxsplit_nw_switch_bb_s0 muxsplit_nw_switch_bb_sl muxsplit_nw_switch_bb_sr vssd0
+ vssio vddio vccd0 vref_w/vddio_q vddio vccd0 w_4981_990174# w_11281_990174# vdda0
+ vssa0 vcap_w/cneg sky130_fd_io__top_amuxsplitv2
Xvdda1_0_pad vref_w/vddio_q vcap_w/cneg vssio vdda1_0 vref_e/amuxbus_b vref_e/amuxbus_a
+ vdda1 vssd0 vccd0 vssa1 vddio vddio vccd0 sky130_ef_io__vdda_hvc_clamped_pad
Xgpio0_1_pad gpio0_1_dm[0] gpio0_1_ib_mode_sel gpio0_1_enable_h gpio0_1_enable_inp_h
+ gpio0_1_slow gpio0_1_vtrip_sel gpio0_1_enable_vddio gpio0_1_enable_vdda_h gpio0_1_pad_a_noesd_h
+ gpio0_1_analog_pol gpio0_1_hld_h_n w_694469_99069# gpio0_1_dm[1] w_692355_95752#
+ gpio0_1_dm[2] w_692253_99070# gpio0_1_pad_a_esd_1_h gpio0_1_tie_hi_esd gpio0_1_enable_vswitch_h
+ gpio0_1_tie_lo_esd gpio0_1_oe_n w_694469_95752# vref_e/amuxbus_b gpio0_1_analog_sel
+ vddio vref_e/amuxbus_a gpio0_1_in_h vddio gpio0_1_inp_dis gpio0_1_out gpio0_1_hld_ovr
+ vccd0 gpio0_1 vccd0 gpio0_1_pad_a_esd_0_h gpio0_1_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio0_1_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio2_4_pad gpio2_4_dm[0] gpio2_4_ib_mode_sel gpio2_4_enable_h gpio2_4_enable_inp_h
+ gpio2_4_slow gpio2_4_vtrip_sel gpio2_4_enable_vddio gpio2_4_enable_vdda_h gpio2_4_pad_a_noesd_h
+ gpio2_4_analog_pol gpio2_4_hld_h_n w_694469_866669# gpio2_4_dm[1] w_692355_863352#
+ gpio2_4_dm[2] w_692253_866670# gpio2_4_pad_a_esd_1_h gpio2_4_tie_hi_esd gpio2_4_enable_vswitch_h
+ gpio2_4_tie_lo_esd gpio2_4_oe_n w_694469_863352# vref_e/amuxbus_b gpio2_4_analog_sel
+ vddio vref_e/amuxbus_a gpio2_4_in_h vddio gpio2_4_inp_dis gpio2_4_out gpio2_4_hld_ovr
+ vccd0 gpio2_4 vccd0 gpio2_4_pad_a_esd_0_h gpio2_4_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio2_4_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio4_7_pad gpio4_7_dm[0] gpio4_7_ib_mode_sel gpio4_7_enable_h gpio4_7_enable_inp_h
+ gpio4_7_slow gpio4_7_vtrip_sel gpio4_7_enable_vddio gpio4_7_enable_vdda_h gpio4_7_pad_a_noesd_h
+ gpio4_7_analog_pol gpio4_7_hld_h_n w_77474_1014469# gpio4_7_dm[1] w_80565_1012355#
+ gpio4_7_dm[2] w_77474_1012253# gpio4_7_pad_a_esd_1_h gpio4_7_tie_hi_esd gpio4_7_enable_vswitch_h
+ gpio4_7_tie_lo_esd gpio4_7_oe_n w_80565_1014469# amuxbus_b_n gpio4_7_analog_sel
+ vddio amuxbus_a_n gpio4_7_in_h vddio gpio4_7_inp_dis gpio4_7_out gpio4_7_hld_ovr
+ vccd0 gpio4_7 vccd0 gpio4_7_pad_a_esd_0_h gpio4_7_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio4_7_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio8_0_pad gpio8_0_dm[0] gpio8_0_ib_mode_sel gpio8_0_enable_h gpio8_0_enable_inp_h
+ gpio8_0_slow gpio8_0_vtrip_sel gpio8_0_enable_vddio gpio8_0_enable_vdda_h gpio8_0_pad_a_noesd_h
+ gpio8_0_analog_pol gpio8_0_hld_h_n w_117469_21253# gpio8_0_dm[1] w_114152_23367#
+ gpio8_0_dm[2] w_117469_23367# gpio8_0_pad_a_esd_1_h gpio8_0_tie_hi_esd gpio8_0_enable_vswitch_h
+ gpio8_0_tie_lo_esd gpio8_0_oe_n w_114152_21253# sio_amuxbus_b gpio8_0_analog_sel
+ vddio sio_amuxbus_a gpio8_0_in_h vddio gpio8_0_inp_dis gpio8_0_out gpio8_0_hld_ovr
+ vccd0 gpio8_0 vccd0 gpio8_0_pad_a_esd_0_h gpio8_0_analog_en vssio vdda3 vref_w/vddio_q
+ vcap_w/cneg vssa3 gpio8_0_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio1_2_connects gpio1_2_one gpio1_2_zero gpio1_2_enable_h gpio1_2_tie_hi_esd gpio1_0_vinref
+ gpio1_2_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xvdda0_0_pad vref_w/vddio_q vcap_w/cneg vssio vdda0_0 amuxbus_b_n amuxbus_a_n vdda0
+ vssd0 vccd0 vssa0 vddio vddio vccd0 sky130_ef_io__vdda_hvc_clamped_pad
Xgpio2_5_connects gpio2_5_tie_lo_esd gpio2_5_in gpio2_5_tie_hi_esd gpio2_5_enable_vddio
+ gpio2_5_slow gpio2_5_pad_a_esd_0_h gpio2_5_pad_a_esd_1_h gpio2_5_dm[1] gpio2_5_pad_a_noesd_h
+ gpio2_5_analog_en gpio2_5_dm[0] gpio2_5_analog_pol gpio2_5_inp_dis gpio2_5_enable_inp_h
+ gpio2_5_enable_h gpio2_5_hld_h_n gpio2_5_analog_sel gpio2_5_dm[2] gpio2_5_hld_ovr
+ gpio2_5_out gpio2_5_enable_vswitch_h gpio2_5_enable_vdda_h gpio2_5_vtrip_sel gpio2_5_ib_mode_sel
+ gpio2_5_oe_n gpio2_5_in_h gpio2_5_one gpio2_5_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio1_4_pad vcap_w/cneg vddio vssio vssd0 vssa1 vref_w/vddio_q vddio vdda1 vccd0
+ vccd0 gpio1_4 vref_e/amuxbus_a vref_e/amuxbus_b gpio1_4_dm[0] gpio1_4_dm[1] gpio1_4_dm[2]
+ gpio1_4_inp_dis gpio1_4_vtrip_sel gpio1_4_ib_mode_sel[0] gpio1_4_ib_mode_sel[1]
+ gpio1_4_slew_ctl[0] gpio1_4_slew_ctl[1] gpio1_4_hys_trim gpio1_4_hld_ovr gpio1_4_enable_h
+ gpio1_4_hld_h_n gpio1_4_enable_vdda_h gpio1_4_analog_en gpio1_4_enable_inp_h gpio1_4_in
+ gpio1_4_in_h vcap_e_cpos gpio1_4_out gpio1_4_analog_pol gpio1_4_analog_sel gpio1_4_slow
+ gpio1_4_oe_n gpio1_4_tie_hi_esd gpio1_4_tie_lo_esd gpio1_4_pad_a_esd_0_h gpio1_4_pad_a_esd_1_h
+ gpio1_4_pad_a_noesd_h gpio1_4_enable_vswitch_h gpio1_4_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xgpio4_1_connects gpio4_1_tie_lo_esd gpio4_1_pad_a_esd_1_h gpio4_1_dm[1] gpio4_1_dm[0]
+ gpio4_1_analog_pol gpio4_1_inp_dis gpio4_1_enable_h gpio4_1_hld_h_n gpio4_1_dm[2]
+ gpio4_1_hld_ovr gpio4_1_out gpio4_1_enable_vswitch_h gpio4_1_enable_vdda_h gpio4_1_vtrip_sel
+ gpio4_1_oe_n gpio4_1_tie_hi_esd gpio4_1_in gpio4_1_enable_vddio gpio4_1_slow gpio4_1_pad_a_esd_0_h
+ gpio4_1_pad_a_noesd_h gpio4_1_analog_en gpio4_1_analog_sel gpio4_1_ib_mode_sel gpio4_1_in_h
+ gpio4_1_zero gpio4_1_one gpio4_1_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio3_7_pad gpio3_7_dm[0] gpio3_7_ib_mode_sel gpio3_7_enable_h gpio3_7_enable_inp_h
+ gpio3_7_slow gpio3_7_vtrip_sel gpio3_7_enable_vddio gpio3_7_enable_vdda_h gpio3_7_pad_a_noesd_h
+ gpio3_7_analog_pol gpio3_7_hld_h_n w_430474_1014469# gpio3_7_dm[1] w_433565_1012355#
+ gpio3_7_dm[2] w_430474_1012253# gpio3_7_pad_a_esd_1_h gpio3_7_tie_hi_esd gpio3_7_enable_vswitch_h
+ gpio3_7_tie_lo_esd gpio3_7_oe_n w_433565_1014469# amuxbus_b_n gpio3_7_analog_sel
+ vddio amuxbus_a_n gpio3_7_in_h vddio gpio3_7_inp_dis gpio3_7_out gpio3_7_hld_ovr
+ vccd0 gpio3_7 vccd0 gpio3_7_pad_a_esd_0_h gpio3_7_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio3_7_in vssd0 sky130_ef_io__gpiov2_pad
Xvssio_6_pad vdda2 vssd0 vssa2 vref_w/amuxbus_a vref_w/amuxbus_b vssio_6 vref_w/vddio_q
+ vddio vssio vddio vcap_w/cneg vccd0 vccd0 sky130_ef_io__vssio_hvc_clamped_pad
Xvccd2_0_pad vdda0 vccd0 vssd2[1] vddio amuxbus_b_n vddio vssio amuxbus_a_n vccd0
+ vccd2_0 vccd2[1] vssd0 vssa0 vref_w/vddio_q vcap_w/cneg sky130_ef_io__vccd_lvc_clamped3_pad
Xselect_connects select_tie_lo_esd select_pad_a_esd_1_h select_dm[1] select_dm[0]
+ select_analog_pol select_inp_dis select_enable_h select_hld_h_n select_dm[2] select_hld_ovr
+ select_out select_enable_vswitch_h select_enable_vdda_h select_vtrip_sel select_oe_n
+ select_tie_hi_esd select_in select_enable_vddio select_slow select_pad_a_esd_0_h
+ select_pad_a_noesd_h select_analog_en select_analog_sel select_ib_mode_sel select_in_h
+ select_zero select_one select_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio7_0_pad gpio7_0_dm[0] gpio7_0_ib_mode_sel gpio7_0_enable_h gpio7_0_enable_inp_h
+ gpio7_0_slow gpio7_0_vtrip_sel gpio7_0_enable_vddio gpio7_0_enable_vdda_h gpio7_0_pad_a_noesd_h
+ gpio7_0_analog_pol gpio7_0_hld_h_n w_21151_275074# gpio7_0_dm[1] w_23367_278165#
+ gpio7_0_dm[2] w_23367_275074# gpio7_0_pad_a_esd_1_h gpio7_0_tie_hi_esd gpio7_0_enable_vswitch_h
+ gpio7_0_tie_lo_esd gpio7_0_oe_n w_21253_278165# vref_w/amuxbus_b gpio7_0_analog_sel
+ vddio vref_w/amuxbus_a gpio7_0_in_h vddio gpio7_0_inp_dis gpio7_0_out gpio7_0_hld_ovr
+ vccd0 gpio7_0 vccd0 gpio7_0_pad_a_esd_0_h gpio7_0_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio7_0_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio5_4_connects gpio5_4_tie_lo_esd gpio5_4_in gpio5_4_tie_hi_esd gpio5_4_enable_vddio
+ gpio5_4_slow gpio5_4_pad_a_esd_0_h gpio5_4_pad_a_esd_1_h gpio5_4_dm[1] gpio5_4_pad_a_noesd_h
+ gpio5_4_analog_en gpio5_4_dm[0] gpio5_4_analog_pol gpio5_4_inp_dis gpio5_4_enable_inp_h
+ gpio5_4_enable_h gpio5_4_hld_h_n gpio5_4_analog_sel gpio5_4_dm[2] gpio5_4_hld_ovr
+ gpio5_4_out gpio5_4_enable_vswitch_h gpio5_4_enable_vdda_h gpio5_4_vtrip_sel gpio5_4_ib_mode_sel
+ gpio5_4_oe_n gpio5_4_in_h gpio5_4_one gpio5_4_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xvddio_7_pad vdda2 vcap_w/cneg vddio vref_w/vddio_q vssd0 vddio_7 vssa2 vref_w/amuxbus_b
+ vref_w/amuxbus_a vddio vccd0 vssio vccd0 sky130_ef_io__vddio_hvc_clamped_pad
Xgpio6_7_connects gpio6_7_one gpio6_7_zero gpio6_7_enable_h gpio6_7_tie_hi_esd gpio6_7_vinref
+ gpio6_7_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xgpio7_0_connects gpio7_0_tie_lo_esd gpio7_0_in gpio7_0_tie_hi_esd gpio7_0_enable_vddio
+ gpio7_0_slow gpio7_0_pad_a_esd_0_h gpio7_0_pad_a_esd_1_h gpio7_0_dm[1] gpio7_0_pad_a_noesd_h
+ gpio7_0_analog_en gpio7_0_dm[0] gpio7_0_analog_pol gpio7_0_inp_dis gpio7_0_enable_inp_h
+ gpio7_0_enable_h gpio7_0_hld_h_n gpio7_0_analog_sel gpio7_0_dm[2] gpio7_0_hld_ovr
+ gpio7_0_out gpio7_0_enable_vswitch_h gpio7_0_enable_vdda_h gpio7_0_vtrip_sel gpio7_0_ib_mode_sel
+ gpio7_0_oe_n gpio7_0_in_h gpio7_0_one gpio7_0_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio0_4_pad gpio0_4_dm[0] gpio0_4_ib_mode_sel gpio0_4_enable_h gpio0_4_enable_inp_h
+ gpio0_4_slow gpio0_4_vtrip_sel gpio0_4_enable_vddio gpio0_4_enable_vdda_h gpio0_4_pad_a_noesd_h
+ gpio0_4_analog_pol gpio0_4_hld_h_n w_694469_202069# gpio0_4_dm[1] w_692355_198752#
+ gpio0_4_dm[2] w_692253_202070# gpio0_4_pad_a_esd_1_h gpio0_4_tie_hi_esd gpio0_4_enable_vswitch_h
+ gpio0_4_tie_lo_esd gpio0_4_oe_n w_694469_198752# vref_e/amuxbus_b gpio0_4_analog_sel
+ vddio vref_e/amuxbus_a gpio0_4_in_h vddio gpio0_4_inp_dis gpio0_4_out gpio0_4_hld_ovr
+ vccd0 gpio0_4 vccd0 gpio0_4_pad_a_esd_0_h gpio0_4_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio0_4_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio2_7_pad gpio2_7_dm[0] gpio2_7_ib_mode_sel gpio2_7_enable_h gpio2_7_enable_inp_h
+ gpio2_7_slow gpio2_7_vtrip_sel gpio2_7_enable_vddio gpio2_7_enable_vdda_h gpio2_7_pad_a_noesd_h
+ gpio2_7_analog_pol gpio2_7_hld_h_n w_694469_929669# gpio2_7_dm[1] w_692355_926352#
+ gpio2_7_dm[2] w_692253_929670# gpio2_7_pad_a_esd_1_h gpio2_7_tie_hi_esd gpio2_7_enable_vswitch_h
+ gpio2_7_tie_lo_esd gpio2_7_oe_n w_694469_926352# vref_e/amuxbus_b gpio2_7_analog_sel
+ vddio vref_e/amuxbus_a gpio2_7_in_h vddio gpio2_7_inp_dis gpio2_7_out gpio2_7_hld_ovr
+ vccd0 gpio2_7 vccd0 gpio2_7_pad_a_esd_0_h gpio2_7_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio2_7_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio8_3_connects gpio8_3_tie_lo_esd gpio8_3_pad_a_esd_1_h gpio8_3_dm[1] gpio8_3_dm[0]
+ gpio8_3_analog_pol gpio8_3_inp_dis gpio8_3_enable_h gpio8_3_hld_h_n gpio8_3_dm[2]
+ gpio8_3_hld_ovr gpio8_3_out gpio8_3_enable_vswitch_h gpio8_3_enable_vdda_h gpio8_3_vtrip_sel
+ gpio8_3_oe_n gpio8_3_tie_hi_esd gpio8_3_in gpio8_3_enable_vddio gpio8_3_slow gpio8_3_pad_a_esd_0_h
+ gpio8_3_pad_a_noesd_h gpio8_3_analog_en gpio8_3_analog_sel gpio8_3_ib_mode_sel gpio8_3_in_h
+ gpio8_3_zero gpio8_3_one gpio8_3_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xvccd1_0_pad vdda1 vccd0 vssd1[1] vddio vref_e/amuxbus_b vddio vssio vref_e/amuxbus_a
+ vccd0 vccd1_0 vccd1[1] vssd0 vssa1 vref_w/vddio_q vcap_w/cneg sky130_ef_io__vccd_lvc_clamped3_pad
Xgpio6_0_pad vcap_w/cneg vddio vssio vssd0 vssa2 vref_w/vddio_q vddio vdda2 vccd0
+ vccd0 gpio6_0 vref_w/amuxbus_a vref_w/amuxbus_b gpio6_0_dm[0] gpio6_0_dm[1] gpio6_0_dm[2]
+ gpio6_0_inp_dis gpio6_0_vtrip_sel gpio6_0_ib_mode_sel[0] gpio6_0_ib_mode_sel[1]
+ gpio6_0_slew_ctl[0] gpio6_0_slew_ctl[1] gpio6_0_hys_trim gpio6_0_hld_ovr gpio6_0_enable_h
+ gpio6_0_hld_h_n gpio6_0_enable_vdda_h gpio6_0_analog_en gpio6_0_enable_inp_h gpio6_0_in
+ gpio6_0_in_h vcap_w_cpos gpio6_0_out gpio6_0_analog_pol gpio6_0_analog_sel gpio6_0_slow
+ gpio6_0_oe_n gpio6_0_tie_hi_esd gpio6_0_tie_lo_esd gpio6_0_pad_a_esd_0_h gpio6_0_pad_a_esd_1_h
+ gpio6_0_pad_a_noesd_h gpio6_0_enable_vswitch_h gpio6_0_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xxo1_pad vccd0 vref_w/vddio_q vccd0 vcap_w/cneg vssd0 sio_amuxbus_b sio_amuxbus_a
+ xo1_core vssa3 vddio vddio vdda3 vssio xo1 sky130_fd_io__top_analog_pad
Xgpio8_3_pad gpio8_3_dm[0] gpio8_3_ib_mode_sel gpio8_3_enable_h gpio8_3_enable_inp_h
+ gpio8_3_slow gpio8_3_vtrip_sel gpio8_3_enable_vddio gpio8_3_enable_vdda_h gpio8_3_pad_a_noesd_h
+ gpio8_3_analog_pol gpio8_3_hld_h_n w_186469_21253# gpio8_3_dm[1] w_183152_23367#
+ gpio8_3_dm[2] w_186469_23367# gpio8_3_pad_a_esd_1_h gpio8_3_tie_hi_esd gpio8_3_enable_vswitch_h
+ gpio8_3_tie_lo_esd gpio8_3_oe_n w_183152_21253# sio_amuxbus_b gpio8_3_analog_sel
+ vddio sio_amuxbus_a gpio8_3_in_h vddio gpio8_3_inp_dis gpio8_3_out gpio8_3_hld_ovr
+ vccd0 gpio8_3 vccd0 gpio8_3_pad_a_esd_0_h gpio8_3_analog_en vssio vdda3 vref_w/vddio_q
+ vcap_w/cneg vssa3 gpio8_3_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio0_2_connects gpio0_2_tie_lo_esd gpio0_2_in gpio0_2_tie_hi_esd gpio0_2_enable_vddio
+ gpio0_2_slow gpio0_2_pad_a_esd_0_h gpio0_2_pad_a_esd_1_h gpio0_2_dm[1] gpio0_2_pad_a_noesd_h
+ gpio0_2_analog_en gpio0_2_dm[0] gpio0_2_analog_pol gpio0_2_inp_dis gpio0_2_enable_inp_h
+ gpio0_2_enable_h gpio0_2_hld_h_n gpio0_2_analog_sel gpio0_2_dm[2] gpio0_2_hld_ovr
+ gpio0_2_out gpio0_2_enable_vswitch_h gpio0_2_enable_vdda_h gpio0_2_vtrip_sel gpio0_2_ib_mode_sel
+ gpio0_2_oe_n gpio0_2_in_h gpio0_2_one gpio0_2_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xvccd0_0_pad vdda3 vccd0 sio_amuxbus_b sio_amuxbus_a vccd0_0 vccd0 vddio vssd0 vssio
+ vssa3 vddio vref_w/vddio_q vcap_w/cneg sky130_ef_io__vccd_lvc_clamped_pad
Xgpio1_7_pad vcap_w/cneg vddio vssio vssd0 vssa1 vref_w/vddio_q vddio vdda1 vccd0
+ vccd0 gpio1_7 vref_e/amuxbus_a vref_e/amuxbus_b gpio1_7_dm[0] gpio1_7_dm[1] gpio1_7_dm[2]
+ gpio1_7_inp_dis gpio1_7_vtrip_sel gpio1_7_ib_mode_sel[0] gpio1_7_ib_mode_sel[1]
+ gpio1_7_slew_ctl[0] gpio1_7_slew_ctl[1] gpio1_7_hys_trim gpio1_7_hld_ovr gpio1_7_enable_h
+ gpio1_7_hld_h_n gpio1_7_enable_vdda_h gpio1_7_analog_en gpio1_7_enable_inp_h gpio1_7_in
+ gpio1_7_in_h vcap_e_cpos gpio1_7_out gpio1_7_analog_pol gpio1_7_analog_sel gpio1_7_slow
+ gpio1_7_oe_n gpio1_7_tie_hi_esd gpio1_7_tie_lo_esd gpio1_7_pad_a_esd_0_h gpio1_7_pad_a_esd_1_h
+ gpio1_7_pad_a_noesd_h gpio1_7_enable_vswitch_h gpio1_7_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xgpio1_5_connects gpio1_5_one gpio1_5_zero gpio1_5_enable_h gpio1_5_tie_hi_esd vcap_e_cpos
+ gpio1_5_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xgpio5_0_pad gpio5_0_dm[0] gpio5_0_ib_mode_sel gpio5_0_enable_h gpio5_0_enable_inp_h
+ gpio5_0_slow gpio5_0_vtrip_sel gpio5_0_enable_vddio gpio5_0_enable_vdda_h gpio5_0_pad_a_noesd_h
+ gpio5_0_analog_pol gpio5_0_hld_h_n w_21151_937674# gpio5_0_dm[1] w_23367_940765#
+ gpio5_0_dm[2] w_23367_937674# gpio5_0_pad_a_esd_1_h gpio5_0_tie_hi_esd gpio5_0_enable_vswitch_h
+ gpio5_0_tie_lo_esd gpio5_0_oe_n w_21253_940765# vref_w/amuxbus_b gpio5_0_analog_sel
+ vddio vref_w/amuxbus_a gpio5_0_in_h vddio gpio5_0_inp_dis gpio5_0_out gpio5_0_hld_ovr
+ vccd0 gpio5_0 vccd0 gpio5_0_pad_a_esd_0_h gpio5_0_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio5_0_in vssd0 sky130_ef_io__gpiov2_pad
Xvssio_9_pad vdda3 vssd0 vssa3 sio_amuxbus_a sio_amuxbus_b vssio_9 vref_w/vddio_q
+ vddio vssio vddio vcap_w/cneg vccd0 vccd0 sky130_ef_io__vssio_hvc_clamped_pad
Xvcap_w vcap_w_cpos vcap_w/cneg vssio vref_w/vddio_q vddio vcap_w/cneg vccd0 vssa2
+ vccd0 vddio vdda2 vssd0 vref_w/amuxbus_b vref_w/amuxbus_a sky130_fd_io__top_vrefcapv2
Xgpio7_3_pad gpio7_3_dm[0] gpio7_3_ib_mode_sel gpio7_3_enable_h gpio7_3_enable_inp_h
+ gpio7_3_slow gpio7_3_vtrip_sel gpio7_3_enable_vddio gpio7_3_enable_vdda_h gpio7_3_pad_a_noesd_h
+ gpio7_3_analog_pol gpio7_3_hld_h_n w_21151_212074# gpio7_3_dm[1] w_23367_215165#
+ gpio7_3_dm[2] w_23367_212074# gpio7_3_pad_a_esd_1_h gpio7_3_tie_hi_esd gpio7_3_enable_vswitch_h
+ gpio7_3_tie_lo_esd gpio7_3_oe_n w_21253_215165# vref_w/amuxbus_b gpio7_3_analog_sel
+ vddio vref_w/amuxbus_a gpio7_3_in_h vddio gpio7_3_inp_dis gpio7_3_out gpio7_3_hld_ovr
+ vccd0 gpio7_3 vccd0 gpio7_3_pad_a_esd_0_h gpio7_3_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio7_3_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio3_1_connects gpio3_1_tie_lo_esd gpio3_1_pad_a_esd_1_h gpio3_1_dm[1] gpio3_1_dm[0]
+ gpio3_1_analog_pol gpio3_1_inp_dis gpio3_1_enable_h gpio3_1_hld_h_n gpio3_1_dm[2]
+ gpio3_1_hld_ovr gpio3_1_out gpio3_1_enable_vswitch_h gpio3_1_enable_vdda_h gpio3_1_vtrip_sel
+ gpio3_1_oe_n gpio3_1_tie_hi_esd gpio3_1_in gpio3_1_enable_vddio gpio3_1_slow gpio3_1_pad_a_esd_0_h
+ gpio3_1_pad_a_noesd_h gpio3_1_analog_en gpio3_1_analog_sel gpio3_1_ib_mode_sel gpio3_1_in_h
+ gpio3_1_zero gpio3_1_one gpio3_1_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio4_4_connects gpio4_4_tie_lo_esd gpio4_4_pad_a_esd_1_h gpio4_4_dm[1] gpio4_4_dm[0]
+ gpio4_4_analog_pol gpio4_4_inp_dis gpio4_4_enable_h gpio4_4_hld_h_n gpio4_4_dm[2]
+ gpio4_4_hld_ovr gpio4_4_out gpio4_4_enable_vswitch_h gpio4_4_enable_vdda_h gpio4_4_vtrip_sel
+ gpio4_4_oe_n gpio4_4_tie_hi_esd gpio4_4_in gpio4_4_enable_vddio gpio4_4_slow gpio4_4_pad_a_esd_0_h
+ gpio4_4_pad_a_noesd_h gpio4_4_analog_en gpio4_4_analog_sel gpio4_4_ib_mode_sel gpio4_4_in_h
+ gpio4_4_zero gpio4_4_one gpio4_4_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio0_7_pad gpio0_7_dm[0] gpio0_7_ib_mode_sel gpio0_7_enable_h gpio0_7_enable_inp_h
+ gpio0_7_slow gpio0_7_vtrip_sel gpio0_7_enable_vddio gpio0_7_enable_vdda_h gpio0_7_pad_a_noesd_h
+ gpio0_7_analog_pol gpio0_7_hld_h_n w_694469_265069# gpio0_7_dm[1] w_692355_261752#
+ gpio0_7_dm[2] w_692253_265070# gpio0_7_pad_a_esd_1_h gpio0_7_tie_hi_esd gpio0_7_enable_vswitch_h
+ gpio0_7_tie_lo_esd gpio0_7_oe_n w_694469_261752# vref_e/amuxbus_b gpio0_7_analog_sel
+ vddio vref_e/amuxbus_a gpio0_7_in_h vddio gpio0_7_inp_dis gpio0_7_out gpio0_7_hld_ovr
+ vccd0 gpio0_7 vccd0 gpio0_7_pad_a_esd_0_h gpio0_7_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio0_7_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio4_0_pad gpio4_0_dm[0] gpio4_0_ib_mode_sel gpio4_0_enable_h gpio4_0_enable_inp_h
+ gpio4_0_slow gpio4_0_vtrip_sel gpio4_0_enable_vddio gpio4_0_enable_vdda_h gpio4_0_pad_a_noesd_h
+ gpio4_0_analog_pol gpio4_0_hld_h_n w_291474_1014469# gpio4_0_dm[1] w_294565_1012355#
+ gpio4_0_dm[2] w_291474_1012253# gpio4_0_pad_a_esd_1_h gpio4_0_tie_hi_esd gpio4_0_enable_vswitch_h
+ gpio4_0_tie_lo_esd gpio4_0_oe_n w_294565_1014469# amuxbus_b_n gpio4_0_analog_sel
+ vddio amuxbus_a_n gpio4_0_in_h vddio gpio4_0_inp_dis gpio4_0_out gpio4_0_hld_ovr
+ vccd0 gpio4_0 vccd0 gpio4_0_pad_a_esd_0_h gpio4_0_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio4_0_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio5_7_connects gpio5_7_tie_lo_esd gpio5_7_in gpio5_7_tie_hi_esd gpio5_7_enable_vddio
+ gpio5_7_slow gpio5_7_pad_a_esd_0_h gpio5_7_pad_a_esd_1_h gpio5_7_dm[1] gpio5_7_pad_a_noesd_h
+ gpio5_7_analog_en gpio5_7_dm[0] gpio5_7_analog_pol gpio5_7_inp_dis gpio5_7_enable_inp_h
+ gpio5_7_enable_h gpio5_7_hld_h_n gpio5_7_analog_sel gpio5_7_dm[2] gpio5_7_hld_ovr
+ gpio5_7_out gpio5_7_enable_vswitch_h gpio5_7_enable_vdda_h gpio5_7_vtrip_sel gpio5_7_ib_mode_sel
+ gpio5_7_oe_n gpio5_7_in_h gpio5_7_one gpio5_7_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio6_0_connects gpio6_0_one gpio6_0_zero gpio6_0_enable_h gpio6_0_tie_hi_esd vcap_w_cpos
+ gpio6_0_tie_lo_esd vccd0 vssd0 chip_io_ovt_connects_horiz
Xvssd2_0_pad vdda0 vcap_w/cneg vssd2[0] vccd0 vssd0 vssa0 amuxbus_b_n amuxbus_a_n
+ vssd2_0 vddio vddio vccd0 vref_w/vddio_q vssio vccd2[0] sky130_ef_io__vssd_lvc_clamped3_pad
Xgpio6_3_pad vcap_w/cneg vddio vssio vssd0 vssa2 vref_w/vddio_q vddio vdda2 vccd0
+ vccd0 gpio6_3 vref_w/amuxbus_a vref_w/amuxbus_b gpio6_3_dm[0] gpio6_3_dm[1] gpio6_3_dm[2]
+ gpio6_3_inp_dis gpio6_3_vtrip_sel gpio6_3_ib_mode_sel[0] gpio6_3_ib_mode_sel[1]
+ gpio6_3_slew_ctl[0] gpio6_3_slew_ctl[1] gpio6_3_hys_trim gpio6_3_hld_ovr gpio6_3_enable_h
+ gpio6_3_hld_h_n gpio6_3_enable_vdda_h gpio6_3_analog_en gpio6_3_enable_inp_h gpio6_3_in
+ gpio6_3_in_h vcap_w_cpos gpio6_3_out gpio6_3_analog_pol gpio6_3_analog_sel gpio6_3_slow
+ gpio6_3_oe_n gpio6_3_tie_hi_esd gpio6_3_tie_lo_esd gpio6_3_pad_a_esd_0_h gpio6_3_pad_a_esd_1_h
+ gpio6_3_pad_a_noesd_h gpio6_3_enable_vswitch_h gpio6_3_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xgpio7_3_connects gpio7_3_tie_lo_esd gpio7_3_in gpio7_3_tie_hi_esd gpio7_3_enable_vddio
+ gpio7_3_slow gpio7_3_pad_a_esd_0_h gpio7_3_pad_a_esd_1_h gpio7_3_dm[1] gpio7_3_pad_a_noesd_h
+ gpio7_3_analog_en gpio7_3_dm[0] gpio7_3_analog_pol gpio7_3_inp_dis gpio7_3_enable_inp_h
+ gpio7_3_enable_h gpio7_3_hld_h_n gpio7_3_analog_sel gpio7_3_dm[2] gpio7_3_hld_ovr
+ gpio7_3_out gpio7_3_enable_vswitch_h gpio7_3_enable_vdda_h gpio7_3_vtrip_sel gpio7_3_ib_mode_sel
+ gpio7_3_oe_n gpio7_3_in_h gpio7_3_one gpio7_3_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio8_6_pad gpio8_6_dm[0] gpio8_6_ib_mode_sel gpio8_6_enable_h gpio8_6_enable_inp_h
+ gpio8_6_slow gpio8_6_vtrip_sel gpio8_6_enable_vddio gpio8_6_enable_vdda_h gpio8_6_pad_a_noesd_h
+ gpio8_6_analog_pol gpio8_6_hld_h_n w_435469_21253# gpio8_6_dm[1] w_432152_23367#
+ gpio8_6_dm[2] w_435469_23367# gpio8_6_pad_a_esd_1_h gpio8_6_tie_hi_esd gpio8_6_enable_vswitch_h
+ gpio8_6_tie_lo_esd gpio8_6_oe_n w_432152_21253# sio_amuxbus_b gpio8_6_analog_sel
+ vddio sio_amuxbus_a gpio8_6_in_h vddio gpio8_6_inp_dis gpio8_6_out gpio8_6_hld_ovr
+ vccd0 gpio8_6 vccd0 gpio8_6_pad_a_esd_0_h gpio8_6_analog_en vssio vdda3 vref_w/vddio_q
+ vcap_w/cneg vssa3 gpio8_6_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio8_6_connects gpio8_6_tie_lo_esd gpio8_6_pad_a_esd_1_h gpio8_6_dm[1] gpio8_6_dm[0]
+ gpio8_6_analog_pol gpio8_6_inp_dis gpio8_6_enable_h gpio8_6_hld_h_n gpio8_6_dm[2]
+ gpio8_6_hld_ovr gpio8_6_out gpio8_6_enable_vswitch_h gpio8_6_enable_vdda_h gpio8_6_vtrip_sel
+ gpio8_6_oe_n gpio8_6_tie_hi_esd gpio8_6_in gpio8_6_enable_vddio gpio8_6_slow gpio8_6_pad_a_esd_0_h
+ gpio8_6_pad_a_noesd_h gpio8_6_analog_en gpio8_6_analog_sel gpio8_6_ib_mode_sel gpio8_6_in_h
+ gpio8_6_zero gpio8_6_one gpio8_6_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio3_0_pad gpio3_0_dm[0] gpio3_0_ib_mode_sel gpio3_0_enable_h gpio3_0_enable_inp_h
+ gpio3_0_slow gpio3_0_vtrip_sel gpio3_0_enable_vddio gpio3_0_enable_vdda_h gpio3_0_pad_a_noesd_h
+ gpio3_0_analog_pol gpio3_0_hld_h_n w_644474_1014469# gpio3_0_dm[1] w_647565_1012355#
+ gpio3_0_dm[2] w_644474_1012253# gpio3_0_pad_a_esd_1_h gpio3_0_tie_hi_esd gpio3_0_enable_vswitch_h
+ gpio3_0_tie_lo_esd gpio3_0_oe_n w_647565_1014469# amuxbus_b_n gpio3_0_analog_sel
+ vddio amuxbus_a_n gpio3_0_in_h vddio gpio3_0_inp_dis gpio3_0_out gpio3_0_hld_ovr
+ vccd0 gpio3_0 vccd0 gpio3_0_pad_a_esd_0_h gpio3_0_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio3_0_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio5_3_pad gpio5_3_dm[0] gpio5_3_ib_mode_sel gpio5_3_enable_h gpio5_3_enable_inp_h
+ gpio5_3_slow gpio5_3_vtrip_sel gpio5_3_enable_vddio gpio5_3_enable_vdda_h gpio5_3_pad_a_noesd_h
+ gpio5_3_analog_pol gpio5_3_hld_h_n w_21151_874674# gpio5_3_dm[1] w_23367_877765#
+ gpio5_3_dm[2] w_23367_874674# gpio5_3_pad_a_esd_1_h gpio5_3_tie_hi_esd gpio5_3_enable_vswitch_h
+ gpio5_3_tie_lo_esd gpio5_3_oe_n w_21253_877765# vref_w/amuxbus_b gpio5_3_analog_sel
+ vddio vref_w/amuxbus_a gpio5_3_in_h vddio gpio5_3_inp_dis gpio5_3_out gpio5_3_hld_ovr
+ vccd0 gpio5_3 vccd0 gpio5_3_pad_a_esd_0_h gpio5_3_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio5_3_in vssd0 sky130_ef_io__gpiov2_pad
Xvssd1_0_pad vdda1 vcap_w/cneg vssd1[0] vccd0 vssd0 vssa1 vref_e/amuxbus_b vref_e/amuxbus_a
+ vssd1_0 vddio vddio vccd0 vref_w/vddio_q vssio vccd1[0] sky130_ef_io__vssd_lvc_clamped3_pad
Xgpio7_6_pad gpio7_6_dm[0] gpio7_6_ib_mode_sel gpio7_6_enable_h gpio7_6_enable_inp_h
+ gpio7_6_slow gpio7_6_vtrip_sel gpio7_6_enable_vddio gpio7_6_enable_vdda_h gpio7_6_pad_a_noesd_h
+ gpio7_6_analog_pol gpio7_6_hld_h_n w_21151_106074# gpio7_6_dm[1] w_23367_109165#
+ gpio7_6_dm[2] w_23367_106074# gpio7_6_pad_a_esd_1_h gpio7_6_tie_hi_esd gpio7_6_enable_vswitch_h
+ gpio7_6_tie_lo_esd gpio7_6_oe_n w_21253_109165# vref_w/amuxbus_b gpio7_6_analog_sel
+ vddio vref_w/amuxbus_a gpio7_6_in_h vddio gpio7_6_inp_dis gpio7_6_out gpio7_6_hld_ovr
+ vccd0 gpio7_6 vccd0 gpio7_6_pad_a_esd_0_h gpio7_6_analog_en vssio vdda2 vref_w/vddio_q
+ vcap_w/cneg vssa2 gpio7_6_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio0_5_connects gpio0_5_tie_lo_esd gpio0_5_in gpio0_5_tie_hi_esd gpio0_5_enable_vddio
+ gpio0_5_slow gpio0_5_pad_a_esd_0_h gpio0_5_pad_a_esd_1_h gpio0_5_dm[1] gpio0_5_pad_a_noesd_h
+ gpio0_5_analog_en gpio0_5_dm[0] gpio0_5_analog_pol gpio0_5_inp_dis gpio0_5_enable_inp_h
+ gpio0_5_enable_h gpio0_5_hld_h_n gpio0_5_analog_sel gpio0_5_dm[2] gpio0_5_hld_ovr
+ gpio0_5_out gpio0_5_enable_vswitch_h gpio0_5_enable_vdda_h gpio0_5_vtrip_sel gpio0_5_ib_mode_sel
+ gpio0_5_oe_n gpio0_5_in_h gpio0_5_one gpio0_5_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xvddio_0_pad vdda1 vcap_w/cneg vddio vref_w/vddio_q vssd0 vddio_0 vssa1 vref_e/amuxbus_b
+ vref_e/amuxbus_a vddio vccd0 vssio vccd0 sky130_ef_io__vddio_hvc_clamped_pad
Xgpio2_1_connects gpio2_1_tie_lo_esd gpio2_1_in gpio2_1_tie_hi_esd gpio2_1_enable_vddio
+ gpio2_1_slow gpio2_1_pad_a_esd_0_h gpio2_1_pad_a_esd_1_h gpio2_1_dm[1] gpio2_1_pad_a_noesd_h
+ gpio2_1_analog_en gpio2_1_dm[0] gpio2_1_analog_pol gpio2_1_inp_dis gpio2_1_enable_inp_h
+ gpio2_1_enable_h gpio2_1_hld_h_n gpio2_1_analog_sel gpio2_1_dm[2] gpio2_1_hld_ovr
+ gpio2_1_out gpio2_1_enable_vswitch_h gpio2_1_enable_vdda_h gpio2_1_vtrip_sel gpio2_1_ib_mode_sel
+ gpio2_1_oe_n gpio2_1_in_h gpio2_1_one gpio2_1_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xgpio2_0_pad gpio2_0_dm[0] gpio2_0_ib_mode_sel gpio2_0_enable_h gpio2_0_enable_inp_h
+ gpio2_0_slow gpio2_0_vtrip_sel gpio2_0_enable_vddio gpio2_0_enable_vdda_h gpio2_0_pad_a_noesd_h
+ gpio2_0_analog_pol gpio2_0_hld_h_n w_694469_762669# gpio2_0_dm[1] w_692355_759352#
+ gpio2_0_dm[2] w_692253_762670# gpio2_0_pad_a_esd_1_h gpio2_0_tie_hi_esd gpio2_0_enable_vswitch_h
+ gpio2_0_tie_lo_esd gpio2_0_oe_n w_694469_759352# vref_e/amuxbus_b gpio2_0_analog_sel
+ vddio vref_e/amuxbus_a gpio2_0_in_h vddio gpio2_0_inp_dis gpio2_0_out gpio2_0_hld_ovr
+ vccd0 gpio2_0 vccd0 gpio2_0_pad_a_esd_0_h gpio2_0_analog_en vssio vdda1 vref_w/vddio_q
+ vcap_w/cneg vssa1 gpio2_0_in vssd0 sky130_ef_io__gpiov2_pad
Xanalog_1_pad vccd0 vref_w/vddio_q vccd0 vcap_w/cneg vssd0 amuxbus_b_n amuxbus_a_n
+ analog_1_core vssa0 vddio vddio vdda0 vssio analog_1 sky130_fd_io__top_analog_pad
Xgpio3_4_connects gpio3_4_tie_lo_esd gpio3_4_pad_a_esd_1_h gpio3_4_dm[1] gpio3_4_dm[0]
+ gpio3_4_analog_pol gpio3_4_inp_dis gpio3_4_enable_h gpio3_4_hld_h_n gpio3_4_dm[2]
+ gpio3_4_hld_ovr gpio3_4_out gpio3_4_enable_vswitch_h gpio3_4_enable_vdda_h gpio3_4_vtrip_sel
+ gpio3_4_oe_n gpio3_4_tie_hi_esd gpio3_4_in gpio3_4_enable_vddio gpio3_4_slow gpio3_4_pad_a_esd_0_h
+ gpio3_4_pad_a_noesd_h gpio3_4_analog_en gpio3_4_analog_sel gpio3_4_ib_mode_sel gpio3_4_in_h
+ gpio3_4_zero gpio3_4_one gpio3_4_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xvssd0_0_pad vdda3 vssd0_0 vccd0 vddio vddio sio_amuxbus_a sio_amuxbus_b vref_w/vddio_q
+ vssd0 vssio vcap_w/cneg vccd0 vssa3 sky130_ef_io__vssd_lvc_clamped_pad
Xgpio4_3_pad gpio4_3_dm[0] gpio4_3_ib_mode_sel gpio4_3_enable_h gpio4_3_enable_inp_h
+ gpio4_3_slow gpio4_3_vtrip_sel gpio4_3_enable_vddio gpio4_3_enable_vdda_h gpio4_3_pad_a_noesd_h
+ gpio4_3_analog_pol gpio4_3_hld_h_n w_219474_1014469# gpio4_3_dm[1] w_222565_1012355#
+ gpio4_3_dm[2] w_219474_1012253# gpio4_3_pad_a_esd_1_h gpio4_3_tie_hi_esd gpio4_3_enable_vswitch_h
+ gpio4_3_tie_lo_esd gpio4_3_oe_n w_222565_1014469# amuxbus_b_n gpio4_3_analog_sel
+ vddio amuxbus_a_n gpio4_3_in_h vddio gpio4_3_inp_dis gpio4_3_out gpio4_3_hld_ovr
+ vccd0 gpio4_3 vccd0 gpio4_3_pad_a_esd_0_h gpio4_3_analog_en vssio vdda0 vref_w/vddio_q
+ vcap_w/cneg vssa0 gpio4_3_in vssd0 sky130_ef_io__gpiov2_pad
Xgpio6_6_pad vcap_w/cneg vddio vssio vssd0 vssa2 vref_w/vddio_q vddio vdda2 vccd0
+ vccd0 gpio6_6 vref_w/amuxbus_a vref_w/amuxbus_b gpio6_6_dm[0] gpio6_6_dm[1] gpio6_6_dm[2]
+ gpio6_6_inp_dis gpio6_6_vtrip_sel gpio6_6_ib_mode_sel[0] gpio6_6_ib_mode_sel[1]
+ gpio6_6_slew_ctl[0] gpio6_6_slew_ctl[1] gpio6_6_hys_trim gpio6_6_hld_ovr gpio6_6_enable_h
+ gpio6_6_hld_h_n gpio6_6_enable_vdda_h gpio6_6_analog_en gpio6_6_enable_inp_h gpio6_6_in
+ gpio6_6_in_h gpio6_7_vinref gpio6_6_out gpio6_6_analog_pol gpio6_6_analog_sel gpio6_6_slow
+ gpio6_6_oe_n gpio6_6_tie_hi_esd gpio6_6_tie_lo_esd gpio6_6_pad_a_esd_0_h gpio6_6_pad_a_esd_1_h
+ gpio6_6_pad_a_noesd_h gpio6_6_enable_vswitch_h gpio6_6_enable_vddio sky130_fd_io__top_gpio_ovtv2
Xgpio4_7_connects gpio4_7_tie_lo_esd gpio4_7_pad_a_esd_1_h gpio4_7_dm[1] gpio4_7_dm[0]
+ gpio4_7_analog_pol gpio4_7_inp_dis gpio4_7_enable_h gpio4_7_hld_h_n gpio4_7_dm[2]
+ gpio4_7_hld_ovr gpio4_7_out gpio4_7_enable_vswitch_h gpio4_7_enable_vdda_h gpio4_7_vtrip_sel
+ gpio4_7_oe_n gpio4_7_tie_hi_esd gpio4_7_in gpio4_7_enable_vddio gpio4_7_slow gpio4_7_pad_a_esd_0_h
+ gpio4_7_pad_a_noesd_h gpio4_7_analog_en gpio4_7_analog_sel gpio4_7_ib_mode_sel gpio4_7_in_h
+ gpio4_7_zero gpio4_7_one gpio4_7_enable_inp_h vccd0 vssd0 chip_io_gpio_connects_vert
Xgpio5_0_connects gpio5_0_tie_lo_esd gpio5_0_in gpio5_0_tie_hi_esd gpio5_0_enable_vddio
+ gpio5_0_slow gpio5_0_pad_a_esd_0_h gpio5_0_pad_a_esd_1_h gpio5_0_dm[1] gpio5_0_pad_a_noesd_h
+ gpio5_0_analog_en gpio5_0_dm[0] gpio5_0_analog_pol gpio5_0_inp_dis gpio5_0_enable_inp_h
+ gpio5_0_enable_h gpio5_0_hld_h_n gpio5_0_analog_sel gpio5_0_dm[2] gpio5_0_hld_ovr
+ gpio5_0_out gpio5_0_enable_vswitch_h gpio5_0_enable_vdda_h gpio5_0_vtrip_sel gpio5_0_ib_mode_sel
+ gpio5_0_oe_n gpio5_0_in_h gpio5_0_one gpio5_0_zero vccd0 vssd0 chip_io_gpio_connects_horiz
Xxi0_pad vccd0 vref_w/vddio_q vccd0 vcap_w/cneg vssd0 sio_amuxbus_b sio_amuxbus_a
+ xi0_core vssa3 vddio vddio vdda3 vssio xi0 sky130_fd_io__top_analog_pad
.ends

