magic
tech sky130A
magscale 1 2
timestamp 1726510233
<< metal1 >>
rect 348 9642 396 16680
rect 346 9636 398 9642
rect 346 9443 398 9449
rect 348 -1482 396 9443
rect 444 -1154 492 16680
rect 540 -792 588 16680
rect 636 911 684 16680
rect 634 905 686 911
rect 634 719 686 726
rect 538 -798 590 -792
rect 538 -856 590 -850
rect 442 -1160 494 -1154
rect 442 -1218 494 -1212
rect 444 -1482 492 -1218
rect 540 -1482 588 -856
rect 636 -1482 684 719
rect 732 279 780 16680
rect 838 4119 845 4411
rect 897 4171 904 4411
rect 897 4119 948 4171
rect 730 273 782 279
rect 730 108 782 114
rect 732 -1482 780 108
<< via1 >>
rect 346 9449 398 9636
rect 634 726 686 905
rect 538 -850 590 -798
rect 442 -1212 494 -1160
rect 845 4119 897 4411
rect 730 114 782 273
<< metal2 >>
rect 0 16572 778 16578
rect 0 16458 655 16572
rect 769 16458 778 16572
rect 0 16454 778 16458
rect 650 16453 778 16454
rect 0 15982 845 15988
rect 0 15936 910 15982
rect 0 15622 401 15674
rect 355 15573 401 15622
rect 355 15527 910 15573
rect 358 15379 910 15431
rect 358 15354 410 15379
rect 0 15302 410 15354
rect 0 14054 910 14106
rect 0 13343 910 13395
rect 0 12134 910 12186
rect 0 11285 910 11337
rect 0 10907 910 10959
rect 0 10556 842 10608
rect 790 10507 842 10556
rect 790 10455 910 10507
rect 0 10242 910 10294
rect 340 9565 346 9636
rect 0 9513 346 9565
rect 340 9449 346 9513
rect 398 9565 404 9636
rect 398 9513 910 9565
rect 398 9449 404 9513
rect 0 8979 526 8983
rect 0 8927 910 8979
rect 0 7556 910 7608
rect 712 7479 786 7484
rect 712 7312 721 7479
rect 0 7263 721 7312
rect 777 7263 786 7479
rect 0 7260 786 7263
rect 712 7258 786 7260
rect 0 6634 910 6686
rect 845 4411 897 4419
rect 0 4346 845 4398
rect 845 4113 897 4119
rect 397 4094 611 4097
rect 0 4088 611 4094
rect 0 3880 402 4088
rect 397 3684 402 3880
rect 606 3684 611 4088
rect 397 3675 611 3684
rect 0 3238 1149 3290
rect 0 2872 910 3002
rect 0 1614 952 1742
rect 0 1314 734 1366
rect 682 1195 734 1314
rect 824 1273 952 1614
rect 682 1143 962 1195
rect 910 1083 962 1143
rect 647 1066 877 1069
rect 0 1064 877 1066
rect 0 1014 656 1064
rect 647 1008 656 1014
rect 867 1008 877 1064
rect 647 1003 877 1008
rect 634 905 910 916
rect 0 726 634 768
rect 686 876 910 905
rect 0 716 686 726
rect 731 808 957 817
rect 731 752 736 808
rect 952 752 957 808
rect 731 743 957 752
rect 731 466 787 743
rect 0 414 787 466
rect 724 166 730 273
rect 0 114 730 166
rect 782 166 788 273
rect 910 166 950 714
rect 782 114 950 166
rect 753 -797 813 -788
rect 0 -850 538 -798
rect 590 -850 753 -798
rect 740 -1017 753 -850
rect 740 -1026 813 -1017
rect 578 -1159 638 -1150
rect 0 -1212 442 -1160
rect 494 -1212 578 -1160
rect 565 -1379 578 -1212
rect 565 -1388 638 -1379
<< via2 >>
rect 655 16458 769 16572
rect 721 7263 777 7479
rect 402 3684 606 4088
rect 656 1008 867 1064
rect 736 752 952 808
rect 753 -1017 813 -797
rect 578 -1379 638 -1159
<< metal3 >>
rect 650 16572 910 16577
rect 650 16458 655 16572
rect 769 16458 910 16572
rect 650 16453 910 16458
rect 716 7479 910 7484
rect 716 7263 721 7479
rect 777 7418 910 7479
rect 777 7263 791 7418
rect 716 7258 791 7263
rect 397 4088 910 4093
rect 397 3684 402 4088
rect 606 3879 910 4088
rect 606 3684 611 3879
rect 397 3675 611 3684
rect 647 1064 877 1069
rect 647 1008 656 1064
rect 867 1008 877 1064
rect 647 1003 877 1008
rect 802 941 877 1003
rect 802 875 910 941
rect 731 808 957 814
rect 731 752 736 808
rect 952 752 957 808
rect 731 743 957 752
rect 2657 17 3616 26
rect 2657 -146 2716 17
rect 3588 -146 3616 17
rect 2657 -154 3616 -146
rect 2657 -484 10158 -474
rect 2657 -647 9258 -484
rect 10130 -647 10158 -484
rect 2657 -654 10158 -647
rect 748 -797 932 -792
rect 748 -1017 753 -797
rect 813 -852 932 -797
rect 813 -1017 818 -852
rect 748 -1022 818 -1017
rect 2657 -983 3616 -974
rect 2657 -1146 2716 -983
rect 3588 -1146 3616 -983
rect 2657 -1154 3616 -1146
rect 573 -1159 643 -1154
rect 573 -1379 578 -1159
rect 638 -1293 643 -1159
rect 638 -1353 935 -1293
rect 638 -1379 643 -1353
rect 573 -1391 643 -1379
rect 2657 -1484 10158 -1474
rect 2657 -1647 9257 -1484
rect 10129 -1647 10158 -1484
rect 2657 -1654 10158 -1647
rect 2657 -1983 3616 -1974
rect 2657 -2146 2716 -1983
rect 3588 -2146 3616 -1983
rect 2657 -2154 3616 -2146
<< via3 >>
rect 2716 -146 3588 17
rect 9258 -647 10130 -484
rect 2716 -1146 3588 -983
rect 9257 -1647 10129 -1484
rect 2716 -2146 3588 -1983
<< metal4 >>
rect 2714 17 3590 19
rect 2714 -146 2716 17
rect 3588 -146 3590 17
rect 2714 -148 3590 -146
rect 9256 -484 10132 -482
rect 9256 -647 9258 -484
rect 10130 -647 10132 -484
rect 9256 -649 10132 -647
rect 2714 -983 3590 -981
rect 2714 -1146 2716 -983
rect 3588 -1146 3590 -983
rect 2714 -1148 3590 -1146
rect 9255 -1484 10131 -1482
rect 9255 -1647 9257 -1484
rect 10129 -1647 10131 -1484
rect 9255 -1649 10131 -1647
rect 2714 -1983 3590 -1981
rect 2714 -2146 2716 -1983
rect 3588 -2146 3590 -1983
rect 2714 -2148 3590 -2146
use constant_block  constant_block_0
timestamp 1706127523
transform 0 -1 3154 -1 0 228
box 146 496 2430 2224
<< labels >>
flabel metal2 s 0 114 200 166 0 FreeSans 320 0 0 0 tie_lo_esd
port 1 nsew
flabel metal2 s 0 2872 200 3002 0 FreeSans 320 0 0 0 pad_a_esd_1_h
port 2 nsew
flabel metal2 s 0 3238 200 3290 0 FreeSans 320 0 0 0 dm[1]
port 3 nsew
flabel metal2 s 0 6634 200 6686 0 FreeSans 320 0 0 0 dm[0]
port 4 nsew
flabel metal2 s 0 7260 200 7312 0 FreeSans 320 0 0 0 analog_pol
port 5 nsew
flabel metal2 s 0 7556 200 7608 0 FreeSans 320 0 0 0 inp_dis
port 6 nsew
flabel metal2 s 0 9513 200 9565 0 FreeSans 320 0 0 0 enable_h
port 7 nsew
flabel metal2 s 0 10242 200 10294 0 FreeSans 320 0 0 0 hld_h_n
port 8 nsew
flabel metal2 s 0 10907 200 10959 0 FreeSans 320 0 0 0 dm[2]
port 9 nsew
flabel metal2 s 0 11285 200 11337 0 FreeSans 320 0 0 0 hld_ovr
port 10 nsew
flabel metal2 s 0 12134 200 12186 0 FreeSans 320 0 0 0 out
port 11 nsew
flabel metal2 s 0 13343 200 13395 0 FreeSans 320 0 0 0 enable_vswitch_h
port 12 nsew
flabel metal2 s 0 14054 200 14106 0 FreeSans 320 0 0 0 enable_vdda_h
port 13 nsew
flabel metal2 s 0 15302 200 15354 0 FreeSans 320 0 0 0 vtrip_sel
port 14 nsew
flabel metal2 s 0 15936 200 15988 0 FreeSans 320 0 0 0 oe_n
port 15 nsew
flabel metal2 s 0 716 200 768 0 FreeSans 320 0 0 0 tie_hi_esd
port 16 nsew
flabel metal2 s 0 414 200 466 0 FreeSans 320 0 0 0 in
port 17 nsew
flabel metal2 s 0 1014 200 1066 0 FreeSans 320 0 0 0 enable_vddio
port 18 nsew
flabel metal2 s 0 1314 200 1366 0 FreeSans 320 0 0 0 slow
port 19 nsew
flabel metal2 s 0 1614 200 1742 0 FreeSans 320 0 0 0 pad_a_esd_0_h
port 20 nsew
flabel metal2 s 0 3880 200 4094 0 FreeSans 320 0 0 0 pad_a_noesd_h
port 21 nsew
flabel metal2 s 0 4346 200 4398 0 FreeSans 320 0 0 0 analog_en
port 22 nsew
flabel metal2 s 0 10556 200 10608 0 FreeSans 320 0 0 0 analog_sel
port 23 nsew
flabel metal2 s 0 15622 200 15674 0 FreeSans 320 0 0 0 ib_mode_sel
port 24 nsew
flabel metal2 s 0 16454 200 16578 0 FreeSans 320 0 0 0 in_h
port 25 nsew
flabel metal2 s 0 8927 200 8983 0 FreeSans 320 0 0 0 enable_inp_h
port 28 nsew
flabel metal2 s 0 -850 200 -798 0 FreeSans 320 0 0 0 zero
port 26 nsew
flabel metal2 s 0 -1212 200 -1160 0 FreeSans 320 0 0 0 one
port 27 nsew
<< properties >>
string FIXED_BBOX 0 657 1317 16656
string flatten true
<< end >>
