magic
tech sky130A
magscale 1 2
timestamp 1706150479
<< checkpaint >>
rect -1074 30142 2013 30165
rect -1074 21312 2056 30142
rect -1074 18554 2066 21312
rect -1074 -3261 2056 18554
rect -1074 -3456 2013 -3261
<< metal2 >>
rect 270 24543 318 28882
rect 266 24534 322 24543
rect 266 24343 322 24354
rect 270 -2001 318 24343
rect 364 -1245 412 28882
rect 458 -793 510 28882
rect 556 2810 604 28882
rect 652 5728 700 28882
rect 748 20052 796 28882
rect 744 20040 800 20052
rect 744 19814 800 19823
rect 640 5712 712 5728
rect 640 5592 648 5712
rect 704 5592 712 5712
rect 640 5575 712 5592
rect 548 2801 613 2810
rect 548 2684 552 2801
rect 608 2684 613 2801
rect 548 2675 613 2684
rect 456 -802 512 -793
rect 456 -1013 512 -1001
rect 359 -1257 415 -1245
rect 359 -1465 415 -1453
rect 364 -2001 412 -1465
rect 458 -2001 510 -1013
rect 556 -2001 604 2675
rect 652 -2001 700 5575
rect 748 -2001 796 19814
<< via2 >>
rect 266 24354 322 24534
rect 744 19823 800 20040
rect 648 5592 704 5712
rect 552 2684 608 2801
rect 456 -1001 512 -802
rect 359 -1453 415 -1257
<< metal3 >>
rect 261 24534 327 24543
rect 261 24354 266 24534
rect 322 24354 327 24534
rect 261 24343 327 24354
rect 738 20040 806 20052
rect 738 19823 744 20040
rect 800 19823 806 20040
rect 738 19814 806 19823
rect 640 5712 712 5728
rect 640 5592 648 5712
rect 704 5592 712 5712
rect 640 5575 712 5592
rect 547 2801 613 2816
rect 547 2684 552 2801
rect 608 2684 613 2801
rect 547 2669 613 2684
rect 2653 -212 3552 -202
rect 2653 -374 2657 -212
rect 3540 -374 3552 -212
rect 2653 -382 3552 -374
rect 2653 -710 10095 -702
rect 451 -802 517 -793
rect 451 -1001 456 -802
rect 512 -1001 517 -802
rect 2653 -876 9167 -710
rect 10079 -876 10095 -710
rect 2653 -882 10095 -876
rect 451 -1032 517 -1001
rect 240 -1102 942 -1032
rect 2653 -1209 3552 -1202
rect 354 -1257 420 -1245
rect 354 -1453 359 -1257
rect 415 -1453 420 -1257
rect 2653 -1371 2657 -1209
rect 3540 -1371 3552 -1209
rect 2653 -1382 3552 -1371
rect 354 -1482 420 -1453
rect 240 -1552 952 -1482
rect 2653 -1709 10095 -1702
rect 2653 -1875 9167 -1709
rect 10079 -1875 10095 -1709
rect 2653 -1882 10095 -1875
rect 2653 -2209 3552 -2202
rect 2653 -2371 2656 -2209
rect 3539 -2371 3552 -2209
rect 2653 -2382 3552 -2371
<< via3 >>
rect 2657 -374 3540 -212
rect 9167 -876 10079 -710
rect 2657 -1371 3540 -1209
rect 9167 -1875 10079 -1709
rect 2656 -2371 3539 -2209
<< metal4 >>
rect 2655 -212 3542 -210
rect 2655 -374 2657 -212
rect 3540 -374 3542 -212
rect 2655 -376 3542 -374
rect 9165 -710 10081 -708
rect 9165 -876 9167 -710
rect 10079 -876 10081 -710
rect 9165 -878 10081 -876
rect 2655 -1209 3542 -1207
rect 2655 -1371 2657 -1209
rect 3540 -1371 3542 -1209
rect 2655 -1373 3542 -1371
rect 9165 -1709 10081 -1707
rect 9165 -1875 9167 -1709
rect 10079 -1875 10081 -1709
rect 9165 -1877 10081 -1875
rect 2654 -2209 3541 -2207
rect 2654 -2371 2656 -2209
rect 3539 -2371 3541 -2209
rect 2654 -2373 3541 -2371
use constant_block  constant_block_0
timestamp 1706127523
transform 0 -1 3149 -1 0 0
box 146 496 2430 2224
<< labels >>
flabel metal3 s 240 -1552 540 -1482 0 FreeSans 320 0 0 0 one
port 27 nsew
flabel metal3 s 240 -1102 540 -1032 0 FreeSans 320 0 0 0 zero
port 28 nsew
<< properties >>
string FIXED_BBOX 240 770 840 28770
string flatten true
<< end >>
