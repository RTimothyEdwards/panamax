magic
tech sky130A
timestamp 1726600844
<< checkpaint >>
rect 258364 19078 261905 19776
rect 258364 17982 262260 19078
rect 259162 13185 262260 17982
<< metal3 >>
rect 261903 19078 262280 19098
rect 261903 18683 261923 19078
rect 262260 18683 262280 19078
rect 261903 18663 262280 18683
rect 259144 18469 259571 18490
rect 259144 18193 259165 18469
rect 259552 18193 259571 18469
rect 259144 18177 259571 18193
rect 260850 18480 261223 18494
rect 260850 18191 260864 18480
rect 261205 18191 261223 18480
rect 260850 18172 261223 18191
rect 260273 16295 260734 16315
rect 260273 16018 260293 16295
rect 260714 16018 260734 16295
rect 260273 15998 260734 16018
rect 261332 15814 261740 15834
rect 261332 15414 261352 15814
rect 261720 15414 261740 15814
rect 261332 15394 261740 15414
rect 260266 14810 260734 14830
rect 260266 14743 260286 14810
rect 260714 14743 260734 14810
rect 260266 14723 260734 14743
rect 259796 13553 260159 13573
rect 259796 13185 259816 13553
rect 260139 13185 260159 13553
rect 259796 13165 260159 13185
<< via3 >>
rect 261923 18683 262260 19078
rect 259165 18193 259552 18469
rect 260864 18191 261205 18480
rect 260293 16018 260714 16295
rect 261352 15414 261720 15814
rect 260286 14743 260714 14810
rect 259816 13185 260139 13553
<< metal4 >>
rect 261903 19078 262280 19098
rect 261903 18683 261923 19078
rect 262260 18683 262280 19078
rect 261903 18663 262280 18683
rect 259144 18469 259571 18490
rect 259144 18193 259165 18469
rect 259552 18193 259571 18469
rect 259144 18177 259571 18193
rect 260850 18480 261223 18494
rect 260850 18191 260864 18480
rect 261205 18191 261223 18480
rect 260850 18172 261223 18191
rect 260273 16295 260734 16315
rect 260273 16018 260293 16295
rect 260714 16018 260734 16295
rect 260273 15998 260734 16018
rect 261332 15814 261740 15834
rect 261332 15414 261352 15814
rect 261720 15414 261740 15814
rect 261332 15394 261740 15414
rect 260266 14810 260734 14830
rect 260266 14743 260286 14810
rect 260714 14743 260734 14810
rect 260266 14723 260734 14743
rect 259796 13553 260159 13573
rect 259796 13185 259816 13553
rect 260139 13185 260159 13553
rect 259796 13165 260159 13185
<< end >>
