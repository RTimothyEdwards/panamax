magic
tech sky130A
timestamp 1746202518
<< fillblock >>
rect 0 0 11269 2202
use font_6C  font_6C_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776550
transform 1 0 2901 0 1 552
box 0 0 180 1260
use font_6E  font_6E_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776997
transform 1 0 3797 0 1 552
box 0 0 540 900
use font_22  font_22_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598785768
transform 1 0 213 0 1 826
box 0 540 540 1260
use font_22  font_22_1
timestamp 1598785768
transform 1 0 10565 0 1 846
box 0 540 540 1260
use font_43  font_43_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763351
transform 1 0 9135 0 1 550
box 0 0 540 1260
use font_49  font_49_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598765816
transform 1 0 8416 0 1 554
box 0 0 540 1260
use font_53  font_53_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768855
transform 1 0 934 0 1 544
box 0 0 540 1260
use font_54  font_54_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768910
transform 1 0 5748 0 1 552
box 0 0 540 1260
use font_61  font_61_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775307
transform 1 0 1652 0 1 548
box 0 0 540 900
use font_65  font_65_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775915
transform 1 0 7179 0 1 546
box 0 0 540 900
use font_67  font_67_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776042
transform 1 0 4517 0 1 552
box 0 -360 540 900
use font_68  font_68_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776130
transform 1 0 6463 0 1 546
box 0 0 540 1260
use font_69  font_69_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776260
transform 1 0 2368 0 1 548
box 0 0 360 1260
use font_69  font_69_1
timestamp 1598776260
transform 1 0 3258 0 1 552
box 0 0 360 1260
use font_73  font_73_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777283
transform 1 0 9853 0 1 544
box 0 0 540 900
<< end >>
