magic
tech sky130A
magscale 1 2
timestamp 1706137558
<< checkpaint >>
rect 26866 5124 31251 6692
rect 23558 3787 31251 5124
rect 13011 3784 31251 3787
rect 10598 3781 31251 3784
rect 10595 1518 31251 3781
rect 7960 -1259 31251 1518
rect 7960 -1414 10878 -1259
rect 12030 -1260 31251 -1259
rect 13011 -1284 31251 -1260
rect 23558 -1820 31251 -1284
rect 26866 -1976 31251 -1820
<< fillblock >>
rect -262 -266 28126 2764
rect -140 -5140 22204 -1424
rect 26 -10348 30014 -6358
use font_2E  font_2E_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598786878
transform 1 0 13290 0 1 0
box 0 0 720 720
use font_4A  font_4A_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598766195
transform 1 0 4704 0 1 -9317
box 0 0 1080 2520
use font_4B  font_4B_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598766293
transform 1 0 20418 0 1 -4282
box 0 0 1080 2520
use font_6B  font_6B_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776472
transform 1 0 1698 0 1 -4282
box 0 0 1080 2520
use font_6C  font_6C_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776550
transform 1 0 8640 0 1 0
box 0 0 360 2520
use font_6C  font_6C_1
timestamp 1598776550
transform 1 0 24780 0 1 -9318
box 0 0 360 2520
use font_6D  font_6D_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776905
transform 1 0 22861 0 1 30
box 0 0 1800 1800
use font_6E  font_6E_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776997
transform 1 0 14658 0 1 -4282
box 0 0 1080 1800
use font_6E  font_6E_1
timestamp 1598776997
transform 1 0 20041 0 1 11
box 0 0 1080 1800
use font_6E  font_6E_2
timestamp 1598776997
transform 1 0 7598 0 1 -9317
box 0 0 1080 1800
use font_6F  font_6F_2 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777049
transform 1 0 10338 0 1 -4282
box 0 0 1080 1800
use font_28  font_28_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1606780629
transform 1 0 250 0 1 -9325
box 0 0 720 2520
use font_29  font_29_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598786350
transform 1 0 2770 0 1 -9325
box 0 0 720 2520
use font_30  font_30_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598786981
transform 1 0 13098 0 1 -9300
box 0 0 1080 2520
use font_30  font_30_1
timestamp 1598786981
transform 1 0 7374 0 1 -4297
box 0 0 1080 2520
use font_30  font_30_2
timestamp 1598786981
transform 1 0 14351 0 1 -7
box 0 0 1080 2520
use font_31  font_31_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787010
transform 1 0 4551 0 1 -4281
box 0 0 1080 2520
use font_32  font_32_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787041
transform 1 0 11658 0 1 -9300
box 0 0 1080 2520
use font_32  font_32_1
timestamp 1598787041
transform 1 0 14538 0 1 -9300
box 0 0 1080 2520
use font_33  font_33_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787077
transform 1 0 5954 0 1 -4297
box 0 0 1080 2520
use font_34  font_34_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787136
transform 1 0 15941 0 1 -9300
box 0 0 1080 2520
use font_37  font_37_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787264
transform 1 0 11855 0 1 1
box 0 0 1080 2520
use font_43  font_43_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763351
transform 1 0 0 0 1 0
box 0 0 1080 2520
use font_43  font_43_1
timestamp 1598763351
transform 1 0 1330 0 1 -9325
box 0 0 1080 2520
use font_44  font_44_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763661
transform 1 0 18978 0 1 -4282
box 0 0 1080 2520
use font_45  font_45_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598765099
transform 1 0 19002 0 1 -9318
box 0 0 1080 2520
use font_50  font_50_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768087
transform 1 0 17538 0 1 -4282
box 0 0 1080 2520
use font_50  font_50_1
timestamp 1598768087
transform 1 0 17171 0 1 7
box 0 0 1080 2520
use font_53  font_53_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768855
transform 1 0 258 0 1 -4282
box 0 0 1080 2520
use font_56  font_56_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598769117
transform 1 0 10455 0 1 15
box 0 0 1080 2520
use font_61  font_61_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775307
transform 1 0 1440 0 1 0
box 0 0 1080 1800
use font_61  font_61_1
timestamp 1598775307
transform 1 0 4320 0 1 0
box 0 0 1080 1800
use font_61  font_61_2
timestamp 1598775307
transform 1 0 21900 0 1 -9318
box 0 0 1080 1800
use font_61  font_61_5
timestamp 1598775307
transform 1 0 18580 0 1 11
box 0 0 1080 1800
use font_61  font_61_6
timestamp 1598775307
transform 1 0 21460 0 1 11
box 0 0 1080 1800
use font_61  font_61_7
timestamp 1598775307
transform 1 0 25000 0 1 11
box 0 0 1080 1800
use font_62  font_62_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775406
transform 1 0 23340 0 1 -9318
box 0 0 1080 2520
use font_65  font_65_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775915
transform 1 0 7200 0 1 0
box 0 0 1080 1800
use font_65  font_65_1
timestamp 1598775915
transform 1 0 9002 0 1 -9334
box 0 0 1080 1800
use font_65  font_65_2
timestamp 1598775915
transform 1 0 25500 0 1 -9318
box 0 0 1080 1800
use font_65  font_65_7
timestamp 1598775915
transform 1 0 13218 0 1 -4282
box 0 0 1080 1800
use font_66  font_66_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775974
transform 1 0 20460 0 1 -9318
box 0 0 1080 2520
use font_70  font_70_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777090
transform 1 0 11778 0 1 -4282
box 0 -720 1080 1800
use font_72  font_72_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777237
transform 1 0 2880 0 1 0
box 0 0 1080 1800
use font_73  font_73_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777283
transform 1 0 26940 0 1 -9318
box 0 0 1080 1800
use font_73  font_73_1
timestamp 1598777283
transform 1 0 28380 0 1 -9318
box 0 0 1080 1800
use font_75  font_75_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777411
transform 1 0 6162 0 1 -9317
box 0 0 1080 1800
use font_76  font_76_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777472
transform 1 0 5760 0 1 0
box 0 0 1080 1800
use font_78  font_78_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777815
transform 1 0 26409 0 1 -24
box 0 0 1080 1800
use font_79  font_79_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777870
transform 1 0 3138 0 1 -4282
box 0 -720 1080 1800
<< end >>
