magic
tech sky130A
magscale 1 2
timestamp 1746115413
<< checkpaint >>
rect 676119 517644 677623 639502
rect 676119 515146 678820 517644
rect 675948 512578 678820 515146
rect 675948 511880 678808 512578
rect 676119 510024 678808 511880
rect 675936 508328 678808 510024
rect 675126 507456 678808 508328
rect 675126 505760 678504 507456
rect 676119 374670 677623 505760
<< metal2 >>
rect 677508 637252 677556 639502
rect 677508 604234 677556 606474
rect 677508 571238 677556 573486
rect 677508 538572 677556 540512
rect 677279 538524 677556 538572
rect 677279 516384 677327 538524
rect 677279 516336 677623 516384
rect 677432 513886 677480 516336
rect 677208 513838 677480 513886
rect 677208 513188 677256 513838
rect 677208 513140 677548 513188
rect 677500 508764 677548 513140
rect 677196 508716 677548 508764
rect 677196 507068 677244 508716
rect 676119 507020 677339 507068
rect 676119 478156 676167 507020
rect 676119 478108 677556 478156
rect 677508 473664 677556 478108
rect 677508 440664 677556 442902
rect 677508 407628 677556 409898
rect 677508 374670 677556 376878
<< properties >>
string flatten true
<< end >>
