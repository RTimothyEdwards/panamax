magic
tech sky130A
magscale 1 2
timestamp 1563081083
<< checkpaint >>
rect 38667 373410 678883 646212
<< metal2 >>
rect 40044 642702 40092 644952
rect 677508 637252 677556 639502
rect 40044 609702 40092 611952
rect 677508 604234 677556 606474
rect 40044 576702 40092 578952
rect 677508 571238 677556 573486
rect 40044 541116 40092 545970
rect 40044 541068 40271 541116
rect 40223 519106 40271 541068
rect 677508 538572 677556 540512
rect 39927 519058 40271 519106
rect 677279 538524 677556 538572
rect 677279 516384 677327 538524
rect 677279 516336 677623 516384
rect 40183 508936 40459 508984
rect 40411 481036 40459 508936
rect 40044 480988 40459 481036
rect 676119 507020 677339 507068
rect 40044 479120 40092 480988
rect 676119 478156 676167 507020
rect 676119 478108 677556 478156
rect 677508 473664 677556 478108
rect 40044 446104 40092 448356
rect 677508 440664 677556 442902
rect 40044 413104 40092 415356
rect 677508 407628 677556 409898
rect 40044 380104 40092 382356
rect 677508 374670 677556 376878
<< end >>
