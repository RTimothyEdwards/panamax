magic
tech sky130A
timestamp 1746204336
<< checkpaint >>
rect -780 5913 2761 6611
rect -780 4817 3116 5913
rect 18 20 3116 4817
<< metal3 >>
rect 2759 5913 3136 5933
rect 2759 5518 2779 5913
rect 3116 5518 3136 5913
rect 2759 5498 3136 5518
rect 0 5304 427 5325
rect 0 5028 21 5304
rect 408 5028 427 5304
rect 0 5012 427 5028
rect 1706 5315 2079 5329
rect 1706 5026 1720 5315
rect 2061 5026 2079 5315
rect 1706 5007 2079 5026
rect 1129 3130 1590 3150
rect 1129 2853 1149 3130
rect 1570 2853 1590 3130
rect 1129 2833 1590 2853
rect 2188 2649 2596 2669
rect 2188 2249 2208 2649
rect 2576 2249 2596 2649
rect 2188 2229 2596 2249
rect 1122 1645 1590 1665
rect 1122 1578 1142 1645
rect 1570 1578 1590 1645
rect 1122 1558 1590 1578
rect 652 388 1015 408
rect 652 20 672 388
rect 995 20 1015 388
rect 652 0 1015 20
<< via3 >>
rect 2779 5518 3116 5913
rect 21 5028 408 5304
rect 1720 5026 2061 5315
rect 1149 2853 1570 3130
rect 2208 2249 2576 2649
rect 1142 1578 1570 1645
rect 672 20 995 388
<< metal4 >>
rect 2759 5913 3136 5933
rect 2759 5518 2779 5913
rect 3116 5518 3136 5913
rect 2759 5498 3136 5518
rect 0 5304 427 5325
rect 0 5028 21 5304
rect 408 5028 427 5304
rect 0 5012 427 5028
rect 1706 5315 2079 5329
rect 1706 5026 1720 5315
rect 2061 5026 2079 5315
rect 1706 5007 2079 5026
rect 1129 3130 1590 3150
rect 1129 2853 1149 3130
rect 1570 2853 1590 3130
rect 1129 2833 1590 2853
rect 2188 2649 2596 2669
rect 2188 2249 2208 2649
rect 2576 2249 2596 2649
rect 2188 2229 2596 2249
rect 1122 1645 1590 1665
rect 1122 1578 1142 1645
rect 1570 1578 1590 1645
rect 1122 1558 1590 1578
rect 652 388 1015 408
rect 652 20 672 388
rect 995 20 1015 388
rect 652 0 1015 20
<< end >>
