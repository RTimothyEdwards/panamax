// Verilog module of padframe panamax generated from layout

`default_nettype none

module panamax (
    `ifdef USE_POWER_PINS
	inout wire	vccd0_0,
	inout wire	vssio_8,
	inout wire	vssd0_0,
	inout wire	vddio_9,
	inout wire	vccd0_1,
	inout wire	vssio_9,
	inout wire	vssa3_0,
	inout wire	vdda3_0,
	inout wire	vssd0_1,
	inout wire	vddio_0,
	inout wire	vssd1_0,
	inout wire	vssio_0,
	inout wire	vddio_1,
	inout wire	vdda1_0,
	inout wire	vssa1_0,
	inout wire	vccd1_0,
	inout wire	vssio_1,
	inout wire	vddio_2,
	inout wire	vdda1_1,
	inout wire	vssa1_1,
	inout wire	vssd1_1,
	inout wire	vssio_2,
	inout wire	vccd1_1,
	inout wire	vddio_3,
	inout wire	vccd2_0,
	inout wire	vssio_4,
	inout wire	vssd2_0,
	inout wire	vssa0_0,
	inout wire	vdda0_0,
	inout wire	vddio_4,
	inout wire	vccd1_2,
	inout wire	vssio_3,
	inout wire	vssd1_2,
	inout wire	vddio_8,
	inout wire	vccd2_2,
	inout wire	vssio_7,
	inout wire	vddio_7,
	inout wire	vdda2_1,
	inout wire	vssa2_1,
	inout wire	vssd2_2,
	inout wire	vssio_6,
	inout wire	vddio_6,
	inout wire	vdda2_0,
	inout wire	vssa2_0,
	inout wire	vccd2_1,
	inout wire	vssio_5,
	inout wire	vssd2_1,
	inout wire	vddio_5,
    `endif /* USE_POWER_PINS */

	inout wire	select,
	input wire	resetb,
	inout wire	gpio8_0,
	inout wire	gpio8_1,
	inout wire	gpio8_2,
	inout wire	gpio8_3,
	inout wire	xi0,
	inout wire	xo0,
	inout wire	xi1,
	inout wire	xo1,
	inout wire	gpio8_4,
	inout wire	gpio8_5,
	inout wire	gpio8_6,
	inout wire	gpio8_7,
	inout wire	sio0,
	inout wire	sio1,
	inout wire	gpio0_0,
	inout wire	gpio0_1,
	inout wire	gpio0_2,
	inout wire	gpio0_3,
	inout wire	gpio0_4,
	inout wire	gpio0_5,
	inout wire	gpio0_6,
	inout wire	gpio0_7,
	inout wire	gpio1_0,
	inout wire	gpio1_1,
	inout wire	gpio1_2,
	inout wire	gpio1_3,
	inout wire	gpio1_4,
	inout wire	gpio1_5,
	inout wire	gpio1_6,
	inout wire	gpio1_7,
	inout wire	gpio2_0,
	inout wire	gpio2_1,
	inout wire	gpio2_2,
	inout wire	gpio2_3,
	inout wire	gpio2_4,
	inout wire	gpio2_5,
	inout wire	gpio2_6,
	inout wire	gpio2_7,
	inout wire	gpio4_7,
	inout wire	gpio4_6,
	inout wire	gpio4_5,
	inout wire	gpio4_4,
	inout wire	gpio4_3,
	inout wire	gpio4_2,
	inout wire	gpio4_1,
	inout wire	gpio4_0,
	inout wire	analog_1,
	inout wire	analog_0,
	inout wire	gpio3_7,
	inout wire	gpio3_6,
	inout wire	gpio3_5,
	inout wire	gpio3_4,
	inout wire	gpio3_3,
	inout wire	gpio3_2,
	inout wire	gpio3_1,
	inout wire	gpio3_0,
	inout wire	gpio7_7,
	inout wire	gpio7_6,
	inout wire	gpio7_5,
	inout wire	gpio7_4,
	inout wire	gpio7_3,
	inout wire	gpio7_2,
	inout wire	gpio7_1,
	inout wire	gpio7_0,
	inout wire	gpio6_7,
	inout wire	gpio6_6,
	inout wire	gpio6_5,
	inout wire	gpio6_4,
	inout wire	gpio6_3,
	inout wire	gpio6_2,
	inout wire	gpio6_1,
	inout wire	gpio6_0,
	inout wire	gpio5_7,
	inout wire	gpio5_6,
	inout wire	gpio5_5,
	inout wire	gpio5_4,
	inout wire	gpio5_3,
	inout wire	gpio5_2,
	inout wire	gpio5_1,
	inout wire	gpio5_0,
	inout wire	vccd0,
	inout wire	vssio,
	inout wire	vssd0,
	inout wire	vddio,
	inout wire	vssa3,
	inout wire	vdda3,
	inout wire	[5:0]	vssd1,
	inout wire	[5:0]	vccd1,
	inout wire	vdda1,
	inout wire	vssa1,
	inout wire	vdda0,
	inout wire	vssa0,
	inout wire	[5:0]	vssd2,
	inout wire	[5:0]	vccd2,
	inout wire	vssa2,
	inout wire	vdda2,
        output wire	[7:0] product_id,
        output wire	[31:0] project_id,
	output wire	select_tie_lo_esd,
	output wire	select_in,
	output wire	select_tie_hi_esd,
	input wire	select_enable_vddio,
	input wire	select_slow,
	inout wire	select_pad_a_esd_0_h,
	inout wire	select_pad_a_esd_1_h,
	inout wire	select_pad_a_noesd_h,
	input wire	select_analog_en,
	input wire	select_analog_pol,
	input wire	select_inp_dis,
	input wire	select_enable_inp_h,
	input wire	select_enable_h,
	input wire	select_hld_h_n,
	input wire	select_analog_sel,
	input wire	[2:0]	select_dm,
	input wire	select_hld_ovr,
	input wire	select_out,
	input wire	select_enable_vswitch_h,
	input wire	select_enable_vdda_h,
	input wire	select_vtrip_sel,
	input wire	select_ib_mode_sel,
	input wire	select_oe_n,
	output wire	select_in_h,
	output wire	select_zero,
	output wire	select_one,
	input wire	resetb_tie_weak_hi_h,
	input wire	resetb_disable_pullup_h,
	output wire	resetb_tie_hi_esd,
	output wire	resetb_xres_h_n,
	output wire	resetb_xres_n,
	output wire	resetb_tie_lo_esd,
	input wire	resetb_inp_sel_h,
	input wire	resetb_en_vddio_sig_h,
	input wire	resetb_filt_in_h,
	inout wire	resetb_pad_a_esd_h,
	input wire	resetb_pullup_h,
	input wire	resetb_enable_h,
	input wire	resetb_enable_vddio,
	output wire	gpio8_0_tie_lo_esd,
	output wire	gpio8_0_in,
	output wire	gpio8_0_tie_hi_esd,
	input wire	gpio8_0_enable_vddio,
	input wire	gpio8_0_slow,
	inout wire	gpio8_0_pad_a_esd_0_h,
	inout wire	gpio8_0_pad_a_esd_1_h,
	inout wire	gpio8_0_pad_a_noesd_h,
	input wire	gpio8_0_analog_en,
	input wire	gpio8_0_analog_pol,
	input wire	gpio8_0_inp_dis,
	input wire	gpio8_0_enable_inp_h,
	input wire	gpio8_0_enable_h,
	input wire	gpio8_0_hld_h_n,
	input wire	gpio8_0_analog_sel,
	input wire	[2:0]	gpio8_0_dm,
	input wire	gpio8_0_hld_ovr,
	input wire	gpio8_0_out,
	input wire	gpio8_0_enable_vswitch_h,
	input wire	gpio8_0_enable_vdda_h,
	input wire	gpio8_0_vtrip_sel,
	input wire	gpio8_0_ib_mode_sel,
	input wire	gpio8_0_oe_n,
	output wire	gpio8_0_in_h,
	output wire	gpio8_0_zero,
	output wire	gpio8_0_one,
	output wire	gpio8_1_tie_lo_esd,
	output wire	gpio8_1_in,
	output wire	gpio8_1_tie_hi_esd,
	input wire	gpio8_1_enable_vddio,
	input wire	gpio8_1_slow,
	inout wire	gpio8_1_pad_a_esd_0_h,
	inout wire	gpio8_1_pad_a_esd_1_h,
	inout wire	gpio8_1_pad_a_noesd_h,
	input wire	gpio8_1_analog_en,
	input wire	gpio8_1_analog_pol,
	input wire	gpio8_1_inp_dis,
	input wire	gpio8_1_enable_inp_h,
	input wire	gpio8_1_enable_h,
	input wire	gpio8_1_hld_h_n,
	input wire	gpio8_1_analog_sel,
	input wire	[2:0]	gpio8_1_dm,
	input wire	gpio8_1_hld_ovr,
	input wire	gpio8_1_out,
	input wire	gpio8_1_enable_vswitch_h,
	input wire	gpio8_1_enable_vdda_h,
	input wire	gpio8_1_vtrip_sel,
	input wire	gpio8_1_ib_mode_sel,
	input wire	gpio8_1_oe_n,
	output wire	gpio8_1_in_h,
	output wire	gpio8_1_zero,
	output wire	gpio8_1_one,
	output wire	gpio8_2_tie_lo_esd,
	output wire	gpio8_2_in,
	output wire	gpio8_2_tie_hi_esd,
	input wire	gpio8_2_enable_vddio,
	input wire	gpio8_2_slow,
	inout wire	gpio8_2_pad_a_esd_0_h,
	inout wire	gpio8_2_pad_a_esd_1_h,
	inout wire	gpio8_2_pad_a_noesd_h,
	input wire	gpio8_2_analog_en,
	input wire	gpio8_2_analog_pol,
	input wire	gpio8_2_inp_dis,
	input wire	gpio8_2_enable_inp_h,
	input wire	gpio8_2_enable_h,
	input wire	gpio8_2_hld_h_n,
	input wire	gpio8_2_analog_sel,
	input wire	[2:0]	gpio8_2_dm,
	input wire	gpio8_2_hld_ovr,
	input wire	gpio8_2_out,
	input wire	gpio8_2_enable_vswitch_h,
	input wire	gpio8_2_enable_vdda_h,
	input wire	gpio8_2_vtrip_sel,
	input wire	gpio8_2_ib_mode_sel,
	input wire	gpio8_2_oe_n,
	output wire	gpio8_2_in_h,
	output wire	gpio8_2_zero,
	output wire	gpio8_2_one,
	output wire	gpio8_3_tie_lo_esd,
	output wire	gpio8_3_in,
	output wire	gpio8_3_tie_hi_esd,
	input wire	gpio8_3_enable_vddio,
	input wire	gpio8_3_slow,
	inout wire	gpio8_3_pad_a_esd_0_h,
	inout wire	gpio8_3_pad_a_esd_1_h,
	inout wire	gpio8_3_pad_a_noesd_h,
	input wire	gpio8_3_analog_en,
	input wire	gpio8_3_analog_pol,
	input wire	gpio8_3_inp_dis,
	input wire	gpio8_3_enable_inp_h,
	input wire	gpio8_3_enable_h,
	input wire	gpio8_3_hld_h_n,
	input wire	gpio8_3_analog_sel,
	input wire	[2:0]	gpio8_3_dm,
	input wire	gpio8_3_hld_ovr,
	input wire	gpio8_3_out,
	input wire	gpio8_3_enable_vswitch_h,
	input wire	gpio8_3_enable_vdda_h,
	input wire	gpio8_3_vtrip_sel,
	input wire	gpio8_3_ib_mode_sel,
	input wire	gpio8_3_oe_n,
	output wire	gpio8_3_in_h,
	output wire	gpio8_3_zero,
	output wire	gpio8_3_one,
	inout wire	xi0_core,
	inout wire	xo0_core,
	inout wire	xi1_core,
	inout wire	xo1_core,
	output wire	gpio8_4_tie_lo_esd,
	output wire	gpio8_4_in,
	output wire	gpio8_4_tie_hi_esd,
	input wire	gpio8_4_enable_vddio,
	input wire	gpio8_4_slow,
	inout wire	gpio8_4_pad_a_esd_0_h,
	inout wire	gpio8_4_pad_a_esd_1_h,
	inout wire	gpio8_4_pad_a_noesd_h,
	input wire	gpio8_4_analog_en,
	input wire	gpio8_4_analog_pol,
	input wire	gpio8_4_inp_dis,
	input wire	gpio8_4_enable_inp_h,
	input wire	gpio8_4_enable_h,
	input wire	gpio8_4_hld_h_n,
	input wire	gpio8_4_analog_sel,
	input wire	[2:0]	gpio8_4_dm,
	input wire	gpio8_4_hld_ovr,
	input wire	gpio8_4_out,
	input wire	gpio8_4_enable_vswitch_h,
	input wire	gpio8_4_enable_vdda_h,
	input wire	gpio8_4_vtrip_sel,
	input wire	gpio8_4_ib_mode_sel,
	input wire	gpio8_4_oe_n,
	output wire	gpio8_4_in_h,
	output wire	gpio8_4_zero,
	output wire	gpio8_4_one,
	output wire	gpio8_5_tie_lo_esd,
	output wire	gpio8_5_in,
	output wire	gpio8_5_tie_hi_esd,
	input wire	gpio8_5_enable_vddio,
	input wire	gpio8_5_slow,
	inout wire	gpio8_5_pad_a_esd_0_h,
	inout wire	gpio8_5_pad_a_esd_1_h,
	inout wire	gpio8_5_pad_a_noesd_h,
	input wire	gpio8_5_analog_en,
	input wire	gpio8_5_analog_pol,
	input wire	gpio8_5_inp_dis,
	input wire	gpio8_5_enable_inp_h,
	input wire	gpio8_5_enable_h,
	input wire	gpio8_5_hld_h_n,
	input wire	gpio8_5_analog_sel,
	input wire	[2:0]	gpio8_5_dm,
	input wire	gpio8_5_hld_ovr,
	input wire	gpio8_5_out,
	input wire	gpio8_5_enable_vswitch_h,
	input wire	gpio8_5_enable_vdda_h,
	input wire	gpio8_5_vtrip_sel,
	input wire	gpio8_5_ib_mode_sel,
	input wire	gpio8_5_oe_n,
	output wire	gpio8_5_in_h,
	output wire	gpio8_5_zero,
	output wire	gpio8_5_one,
	output wire	gpio8_6_tie_lo_esd,
	output wire	gpio8_6_in,
	output wire	gpio8_6_tie_hi_esd,
	input wire	gpio8_6_enable_vddio,
	input wire	gpio8_6_slow,
	inout wire	gpio8_6_pad_a_esd_0_h,
	inout wire	gpio8_6_pad_a_esd_1_h,
	inout wire	gpio8_6_pad_a_noesd_h,
	input wire	gpio8_6_analog_en,
	input wire	gpio8_6_analog_pol,
	input wire	gpio8_6_inp_dis,
	input wire	gpio8_6_enable_inp_h,
	input wire	gpio8_6_enable_h,
	input wire	gpio8_6_hld_h_n,
	input wire	gpio8_6_analog_sel,
	input wire	[2:0]	gpio8_6_dm,
	input wire	gpio8_6_hld_ovr,
	input wire	gpio8_6_out,
	input wire	gpio8_6_enable_vswitch_h,
	input wire	gpio8_6_enable_vdda_h,
	input wire	gpio8_6_vtrip_sel,
	input wire	gpio8_6_ib_mode_sel,
	input wire	gpio8_6_oe_n,
	output wire	gpio8_6_in_h,
	output wire	gpio8_6_zero,
	output wire	gpio8_6_one,
	output wire	gpio8_7_tie_lo_esd,
	output wire	gpio8_7_in,
	output wire	gpio8_7_tie_hi_esd,
	input wire	gpio8_7_enable_vddio,
	input wire	gpio8_7_slow,
	inout wire	gpio8_7_pad_a_esd_0_h,
	inout wire	gpio8_7_pad_a_esd_1_h,
	inout wire	gpio8_7_pad_a_noesd_h,
	input wire	gpio8_7_analog_en,
	input wire	gpio8_7_analog_pol,
	input wire	gpio8_7_inp_dis,
	input wire	gpio8_7_enable_inp_h,
	input wire	gpio8_7_enable_h,
	input wire	gpio8_7_hld_h_n,
	input wire	gpio8_7_analog_sel,
	input wire	[2:0]	gpio8_7_dm,
	input wire	gpio8_7_hld_ovr,
	input wire	gpio8_7_out,
	input wire	gpio8_7_enable_vswitch_h,
	input wire	gpio8_7_enable_vdda_h,
	input wire	gpio8_7_vtrip_sel,
	input wire	gpio8_7_ib_mode_sel,
	input wire	gpio8_7_oe_n,
	output wire	gpio8_7_in_h,
	output wire	gpio8_7_zero,
	output wire	gpio8_7_one,
	output wire	pwrdet_out2_vddio_hv,
	output wire	pwrdet_out1_vddd_hv,
	input wire	pwrdet_in1_vddio_hv,
	input wire	pwrdet_in2_vddd_hv,
	input wire	pwrdet_in1_vddd_hv,
	output wire	pwrdet_out1_vddio_hv,
	output wire	pwrdet_out2_vddd_hv,
	output wire	pwrdet_out3_vddd_hv,
	output wire	pwrdet_vddio_present_vddd_hv,
	output wire	pwrdet_out3_vddio_hv,
	output wire	pwrdet_tie_lo_esd,
	input wire	pwrdet_in3_vddd_hv,
	output wire	pwrdet_vddd_present_vddio_hv,
	input wire	pwrdet_in2_vddio_hv,
	input wire	pwrdet_in3_vddio_hv,
	input wire	pwrdet_rst_por_hv_n,
	inout wire	sio_vinref_dft,
	inout wire	sio_voutref_dft,
	input wire	[1:0]	sio_vref_sel,
	input wire	sio_enable_vdda_h,
	input wire	sio_dft_refgen,
	input wire	[2:0]	sio_voh_sel,
	inout wire	amuxbus_a_n,
	inout wire	amuxbus_b_n,
	inout wire	sio_amuxbus_b,
	inout wire	sio_amuxbus_a,
	input wire	sio_vreg_en_refgen,
	input wire	sio_ibuf_sel_refgen,
	input wire	sio_vohref,
	input wire	sio_hld_h_n_refgen,
	input wire	sio_vtrip_sel_refgen,
	input wire	[1:0]	sio_pad_a_esd_0_h,
	input wire	[1:0]	sio_pad_a_noesd_h,
	input wire	[1:0]	sio_inp_dis,
	output wire	[1:0]	sio_tie_lo_esd,
	input wire	[1:0]	sio_out,
	input wire	[1:0]	sio_vtrip_sel,
	input wire	[1:0]	sio_ibuf_sel,
	input wire	[1:0]	sio_hld_h_n,
	input wire	[1:0]	sio_hld_ovr,
	output wire	[1:0]	sio_in,
	output wire	[1:0]	sio_in_h,
	input wire	[1:0]	sio_oe_n,
	input wire	[1:0]	sio_slow,
	input wire	[1:0]	sio_vreg_en,
	input wire	sio_enable_h,
	input wire	[2:0]	sio_dm1,
	inout wire	[1:0]	sio_pad_a_esd_1_h,
	input wire	[2:0]	sio_dm0,
	input wire	muxsplit_se_hld_vdda_h_n,
	input wire	muxsplit_se_enable_vdda_h,
	input wire	muxsplit_se_switch_aa_sl,
	input wire	muxsplit_se_switch_aa_s0,
	input wire	muxsplit_se_switch_bb_s0,
	input wire	muxsplit_se_switch_bb_sl,
	input wire	muxsplit_se_switch_bb_sr,
	input wire	muxsplit_se_switch_aa_sr,
	output wire	gpio0_0_tie_lo_esd,
	output wire	gpio0_0_in,
	output wire	gpio0_0_tie_hi_esd,
	input wire	gpio0_0_enable_vddio,
	input wire	gpio0_0_slow,
	inout wire	gpio0_0_pad_a_esd_0_h,
	inout wire	gpio0_0_pad_a_esd_1_h,
	inout wire	gpio0_0_pad_a_noesd_h,
	input wire	gpio0_0_analog_en,
	input wire	gpio0_0_analog_pol,
	input wire	gpio0_0_inp_dis,
	input wire	gpio0_0_enable_inp_h,
	input wire	gpio0_0_enable_h,
	input wire	gpio0_0_hld_h_n,
	input wire	gpio0_0_analog_sel,
	input wire	[2:0]	gpio0_0_dm,
	input wire	gpio0_0_hld_ovr,
	input wire	gpio0_0_out,
	input wire	gpio0_0_enable_vswitch_h,
	input wire	gpio0_0_enable_vdda_h,
	input wire	gpio0_0_vtrip_sel,
	input wire	gpio0_0_ib_mode_sel,
	input wire	gpio0_0_oe_n,
	output wire	gpio0_0_in_h,
	output wire	gpio0_0_zero,
	output wire	gpio0_0_one,
	output wire	gpio0_1_tie_lo_esd,
	output wire	gpio0_1_in,
	output wire	gpio0_1_tie_hi_esd,
	input wire	gpio0_1_enable_vddio,
	input wire	gpio0_1_slow,
	inout wire	gpio0_1_pad_a_esd_0_h,
	inout wire	gpio0_1_pad_a_esd_1_h,
	inout wire	gpio0_1_pad_a_noesd_h,
	input wire	gpio0_1_analog_en,
	input wire	gpio0_1_analog_pol,
	input wire	gpio0_1_inp_dis,
	input wire	gpio0_1_enable_inp_h,
	input wire	gpio0_1_enable_h,
	input wire	gpio0_1_hld_h_n,
	input wire	gpio0_1_analog_sel,
	input wire	[2:0]	gpio0_1_dm,
	input wire	gpio0_1_hld_ovr,
	input wire	gpio0_1_out,
	input wire	gpio0_1_enable_vswitch_h,
	input wire	gpio0_1_enable_vdda_h,
	input wire	gpio0_1_vtrip_sel,
	input wire	gpio0_1_ib_mode_sel,
	input wire	gpio0_1_oe_n,
	output wire	gpio0_1_in_h,
	output wire	gpio0_1_zero,
	output wire	gpio0_1_one,
	output wire	gpio0_2_tie_lo_esd,
	output wire	gpio0_2_in,
	output wire	gpio0_2_tie_hi_esd,
	input wire	gpio0_2_enable_vddio,
	input wire	gpio0_2_slow,
	inout wire	gpio0_2_pad_a_esd_0_h,
	inout wire	gpio0_2_pad_a_esd_1_h,
	inout wire	gpio0_2_pad_a_noesd_h,
	input wire	gpio0_2_analog_en,
	input wire	gpio0_2_analog_pol,
	input wire	gpio0_2_inp_dis,
	input wire	gpio0_2_enable_inp_h,
	input wire	gpio0_2_enable_h,
	input wire	gpio0_2_hld_h_n,
	input wire	gpio0_2_analog_sel,
	input wire	[2:0]	gpio0_2_dm,
	input wire	gpio0_2_hld_ovr,
	input wire	gpio0_2_out,
	input wire	gpio0_2_enable_vswitch_h,
	input wire	gpio0_2_enable_vdda_h,
	input wire	gpio0_2_vtrip_sel,
	input wire	gpio0_2_ib_mode_sel,
	input wire	gpio0_2_oe_n,
	output wire	gpio0_2_in_h,
	output wire	gpio0_2_zero,
	output wire	gpio0_2_one,
	output wire	gpio0_3_tie_lo_esd,
	output wire	gpio0_3_in,
	output wire	gpio0_3_tie_hi_esd,
	input wire	gpio0_3_enable_vddio,
	input wire	gpio0_3_slow,
	inout wire	gpio0_3_pad_a_esd_0_h,
	inout wire	gpio0_3_pad_a_esd_1_h,
	inout wire	gpio0_3_pad_a_noesd_h,
	input wire	gpio0_3_analog_en,
	input wire	gpio0_3_analog_pol,
	input wire	gpio0_3_inp_dis,
	input wire	gpio0_3_enable_inp_h,
	input wire	gpio0_3_enable_h,
	input wire	gpio0_3_hld_h_n,
	input wire	gpio0_3_analog_sel,
	input wire	[2:0]	gpio0_3_dm,
	input wire	gpio0_3_hld_ovr,
	input wire	gpio0_3_out,
	input wire	gpio0_3_enable_vswitch_h,
	input wire	gpio0_3_enable_vdda_h,
	input wire	gpio0_3_vtrip_sel,
	input wire	gpio0_3_ib_mode_sel,
	input wire	gpio0_3_oe_n,
	output wire	gpio0_3_in_h,
	output wire	gpio0_3_zero,
	output wire	gpio0_3_one,
	output wire	gpio0_4_tie_lo_esd,
	output wire	gpio0_4_in,
	output wire	gpio0_4_tie_hi_esd,
	input wire	gpio0_4_enable_vddio,
	input wire	gpio0_4_slow,
	inout wire	gpio0_4_pad_a_esd_0_h,
	inout wire	gpio0_4_pad_a_esd_1_h,
	inout wire	gpio0_4_pad_a_noesd_h,
	input wire	gpio0_4_analog_en,
	input wire	gpio0_4_analog_pol,
	input wire	gpio0_4_inp_dis,
	input wire	gpio0_4_enable_inp_h,
	input wire	gpio0_4_enable_h,
	input wire	gpio0_4_hld_h_n,
	input wire	gpio0_4_analog_sel,
	input wire	[2:0]	gpio0_4_dm,
	input wire	gpio0_4_hld_ovr,
	input wire	gpio0_4_out,
	input wire	gpio0_4_enable_vswitch_h,
	input wire	gpio0_4_enable_vdda_h,
	input wire	gpio0_4_vtrip_sel,
	input wire	gpio0_4_ib_mode_sel,
	input wire	gpio0_4_oe_n,
	output wire	gpio0_4_in_h,
	output wire	gpio0_4_zero,
	output wire	gpio0_4_one,
	output wire	gpio0_5_tie_lo_esd,
	output wire	gpio0_5_in,
	output wire	gpio0_5_tie_hi_esd,
	input wire	gpio0_5_enable_vddio,
	input wire	gpio0_5_slow,
	inout wire	gpio0_5_pad_a_esd_0_h,
	inout wire	gpio0_5_pad_a_esd_1_h,
	inout wire	gpio0_5_pad_a_noesd_h,
	input wire	gpio0_5_analog_en,
	input wire	gpio0_5_analog_pol,
	input wire	gpio0_5_inp_dis,
	input wire	gpio0_5_enable_inp_h,
	input wire	gpio0_5_enable_h,
	input wire	gpio0_5_hld_h_n,
	input wire	gpio0_5_analog_sel,
	input wire	[2:0]	gpio0_5_dm,
	input wire	gpio0_5_hld_ovr,
	input wire	gpio0_5_out,
	input wire	gpio0_5_enable_vswitch_h,
	input wire	gpio0_5_enable_vdda_h,
	input wire	gpio0_5_vtrip_sel,
	input wire	gpio0_5_ib_mode_sel,
	input wire	gpio0_5_oe_n,
	output wire	gpio0_5_in_h,
	output wire	gpio0_5_zero,
	output wire	gpio0_5_one,
	output wire	gpio0_6_tie_lo_esd,
	output wire	gpio0_6_in,
	output wire	gpio0_6_tie_hi_esd,
	input wire	gpio0_6_enable_vddio,
	input wire	gpio0_6_slow,
	inout wire	gpio0_6_pad_a_esd_0_h,
	inout wire	gpio0_6_pad_a_esd_1_h,
	inout wire	gpio0_6_pad_a_noesd_h,
	input wire	gpio0_6_analog_en,
	input wire	gpio0_6_analog_pol,
	input wire	gpio0_6_inp_dis,
	input wire	gpio0_6_enable_inp_h,
	input wire	gpio0_6_enable_h,
	input wire	gpio0_6_hld_h_n,
	input wire	gpio0_6_analog_sel,
	input wire	[2:0]	gpio0_6_dm,
	input wire	gpio0_6_hld_ovr,
	input wire	gpio0_6_out,
	input wire	gpio0_6_enable_vswitch_h,
	input wire	gpio0_6_enable_vdda_h,
	input wire	gpio0_6_vtrip_sel,
	input wire	gpio0_6_ib_mode_sel,
	input wire	gpio0_6_oe_n,
	output wire	gpio0_6_in_h,
	output wire	gpio0_6_zero,
	output wire	gpio0_6_one,
	output wire	gpio0_7_tie_lo_esd,
	output wire	gpio0_7_in,
	output wire	gpio0_7_tie_hi_esd,
	input wire	gpio0_7_enable_vddio,
	input wire	gpio0_7_slow,
	inout wire	gpio0_7_pad_a_esd_0_h,
	inout wire	gpio0_7_pad_a_esd_1_h,
	inout wire	gpio0_7_pad_a_noesd_h,
	input wire	gpio0_7_analog_en,
	input wire	gpio0_7_analog_pol,
	input wire	gpio0_7_inp_dis,
	input wire	gpio0_7_enable_inp_h,
	input wire	gpio0_7_enable_h,
	input wire	gpio0_7_hld_h_n,
	input wire	gpio0_7_analog_sel,
	input wire	[2:0]	gpio0_7_dm,
	input wire	gpio0_7_hld_ovr,
	input wire	gpio0_7_out,
	input wire	gpio0_7_enable_vswitch_h,
	input wire	gpio0_7_enable_vdda_h,
	input wire	gpio0_7_vtrip_sel,
	input wire	gpio0_7_ib_mode_sel,
	input wire	gpio0_7_oe_n,
	output wire	gpio0_7_in_h,
	output wire	gpio0_7_zero,
	output wire	gpio0_7_one,
	output wire	gpio1_0_tie_hi_esd,
	input wire	[2:0]	gpio1_0_dm,
	input wire	gpio1_0_slow,
	input wire	gpio1_0_oe_n,
	output wire	gpio1_0_tie_lo_esd,
	input wire	gpio1_0_inp_dis,
	input wire	gpio1_0_enable_vddio,
	input wire	gpio1_0_vtrip_sel,
	input wire	[1:0]	gpio1_0_ib_mode_sel,
	input wire	gpio1_0_out,
	input wire	[1:0]	gpio1_0_slew_ctl,
	input wire	gpio1_0_analog_pol,
	input wire	gpio1_0_analog_sel,
	input wire	gpio1_0_hys_trim,
	input wire	gpio1_0_hld_ovr,
	output wire	gpio1_0_in_h,
	input wire	gpio1_0_enable_h,
	output wire	gpio1_0_in,
	input wire	gpio1_0_hld_h_n,
	input wire	gpio1_0_enable_vdda_h,
	input wire	gpio1_0_analog_en,
	input wire	gpio1_0_enable_inp_h,
	input wire	gpio1_0_enable_vswitch_h,
	inout wire	gpio1_0_pad_a_noesd_h,
	inout wire	gpio1_0_pad_a_esd_0_h,
	inout wire	gpio1_0_pad_a_esd_1_h,
	output wire	gpio1_0_zero,
	output wire	gpio1_0_one,
	output wire	gpio1_1_tie_hi_esd,
	input wire	[2:0]	gpio1_1_dm,
	input wire	gpio1_1_slow,
	input wire	gpio1_1_oe_n,
	output wire	gpio1_1_tie_lo_esd,
	input wire	gpio1_1_inp_dis,
	input wire	gpio1_1_enable_vddio,
	input wire	gpio1_1_vtrip_sel,
	input wire	[1:0]	gpio1_1_ib_mode_sel,
	input wire	gpio1_1_out,
	input wire	[1:0]	gpio1_1_slew_ctl,
	input wire	gpio1_1_analog_pol,
	input wire	gpio1_1_analog_sel,
	input wire	gpio1_1_hys_trim,
	input wire	gpio1_1_hld_ovr,
	output wire	gpio1_1_in_h,
	input wire	gpio1_1_enable_h,
	output wire	gpio1_1_in,
	input wire	gpio1_1_hld_h_n,
	input wire	gpio1_1_enable_vdda_h,
	input wire	gpio1_1_analog_en,
	input wire	gpio1_1_enable_inp_h,
	input wire	gpio1_1_enable_vswitch_h,
	inout wire	gpio1_1_pad_a_noesd_h,
	inout wire	gpio1_1_pad_a_esd_0_h,
	inout wire	gpio1_1_pad_a_esd_1_h,
	output wire	gpio1_1_zero,
	output wire	gpio1_1_one,
	output wire	gpio1_2_tie_hi_esd,
	input wire	[2:0]	gpio1_2_dm,
	input wire	gpio1_2_slow,
	input wire	gpio1_2_oe_n,
	output wire	gpio1_2_tie_lo_esd,
	input wire	gpio1_2_inp_dis,
	input wire	gpio1_2_enable_vddio,
	input wire	gpio1_2_vtrip_sel,
	input wire	[1:0]	gpio1_2_ib_mode_sel,
	input wire	gpio1_2_out,
	input wire	[1:0]	gpio1_2_slew_ctl,
	input wire	gpio1_2_analog_pol,
	input wire	gpio1_2_analog_sel,
	input wire	gpio1_2_hys_trim,
	input wire	gpio1_2_hld_ovr,
	output wire	gpio1_2_in_h,
	input wire	gpio1_2_enable_h,
	output wire	gpio1_2_in,
	input wire	gpio1_2_hld_h_n,
	input wire	gpio1_2_enable_vdda_h,
	input wire	gpio1_2_analog_en,
	input wire	gpio1_2_enable_inp_h,
	input wire	gpio1_2_enable_vswitch_h,
	inout wire	gpio1_2_pad_a_noesd_h,
	inout wire	gpio1_2_pad_a_esd_0_h,
	inout wire	gpio1_2_pad_a_esd_1_h,
	output wire	gpio1_2_zero,
	output wire	gpio1_2_one,
	output wire	gpio1_3_tie_hi_esd,
	input wire	[2:0]	gpio1_3_dm,
	input wire	gpio1_3_slow,
	input wire	gpio1_3_oe_n,
	output wire	gpio1_3_tie_lo_esd,
	input wire	gpio1_3_inp_dis,
	input wire	gpio1_3_enable_vddio,
	input wire	gpio1_3_vtrip_sel,
	input wire	[1:0]	gpio1_3_ib_mode_sel,
	input wire	gpio1_3_out,
	input wire	[1:0]	gpio1_3_slew_ctl,
	input wire	gpio1_3_analog_pol,
	input wire	gpio1_3_analog_sel,
	input wire	gpio1_3_hys_trim,
	input wire	gpio1_3_hld_ovr,
	output wire	gpio1_3_in_h,
	input wire	gpio1_3_enable_h,
	output wire	gpio1_3_in,
	input wire	gpio1_3_hld_h_n,
	input wire	gpio1_3_enable_vdda_h,
	input wire	gpio1_3_analog_en,
	input wire	gpio1_3_enable_inp_h,
	input wire	gpio1_3_enable_vswitch_h,
	inout wire	gpio1_3_pad_a_noesd_h,
	inout wire	gpio1_3_pad_a_esd_0_h,
	inout wire	gpio1_3_pad_a_esd_1_h,
	output wire	gpio1_3_zero,
	output wire	gpio1_3_one,
	input wire	[4:0]	vref_e_ref_sel,
	inout wire	vref_e_vinref,
	input wire	vref_e_enable_h,
	input wire	vref_e_hld_h_n,
	input wire	vref_e_vrefgen_en,
	output wire	gpio1_4_tie_hi_esd,
	input wire	[2:0]	gpio1_4_dm,
	input wire	gpio1_4_slow,
	input wire	gpio1_4_oe_n,
	output wire	gpio1_4_tie_lo_esd,
	input wire	gpio1_4_inp_dis,
	input wire	gpio1_4_enable_vddio,
	input wire	gpio1_4_vtrip_sel,
	input wire	[1:0]	gpio1_4_ib_mode_sel,
	input wire	gpio1_4_out,
	input wire	[1:0]	gpio1_4_slew_ctl,
	input wire	gpio1_4_analog_pol,
	input wire	gpio1_4_analog_sel,
	input wire	gpio1_4_hys_trim,
	input wire	gpio1_4_hld_ovr,
	output wire	gpio1_4_in_h,
	input wire	gpio1_4_enable_h,
	output wire	gpio1_4_in,
	input wire	gpio1_4_hld_h_n,
	input wire	gpio1_4_enable_vdda_h,
	input wire	gpio1_4_analog_en,
	input wire	gpio1_4_enable_inp_h,
	input wire	gpio1_4_enable_vswitch_h,
	inout wire	gpio1_4_pad_a_noesd_h,
	inout wire	gpio1_4_pad_a_esd_0_h,
	inout wire	gpio1_4_pad_a_esd_1_h,
	output wire	gpio1_4_zero,
	output wire	gpio1_4_one,
	output wire	gpio1_5_tie_hi_esd,
	input wire	[2:0]	gpio1_5_dm,
	input wire	gpio1_5_slow,
	input wire	gpio1_5_oe_n,
	output wire	gpio1_5_tie_lo_esd,
	input wire	gpio1_5_inp_dis,
	input wire	gpio1_5_enable_vddio,
	input wire	gpio1_5_vtrip_sel,
	input wire	[1:0]	gpio1_5_ib_mode_sel,
	input wire	gpio1_5_out,
	input wire	[1:0]	gpio1_5_slew_ctl,
	input wire	gpio1_5_analog_pol,
	input wire	gpio1_5_analog_sel,
	input wire	gpio1_5_hys_trim,
	input wire	gpio1_5_hld_ovr,
	output wire	gpio1_5_in_h,
	input wire	gpio1_5_enable_h,
	output wire	gpio1_5_in,
	input wire	gpio1_5_hld_h_n,
	input wire	gpio1_5_enable_vdda_h,
	input wire	gpio1_5_analog_en,
	input wire	gpio1_5_enable_inp_h,
	input wire	gpio1_5_enable_vswitch_h,
	inout wire	gpio1_5_pad_a_noesd_h,
	inout wire	gpio1_5_pad_a_esd_0_h,
	inout wire	gpio1_5_pad_a_esd_1_h,
	output wire	gpio1_5_zero,
	output wire	gpio1_5_one,
	output wire	gpio1_6_tie_hi_esd,
	input wire	[2:0]	gpio1_6_dm,
	input wire	gpio1_6_slow,
	input wire	gpio1_6_oe_n,
	output wire	gpio1_6_tie_lo_esd,
	input wire	gpio1_6_inp_dis,
	input wire	gpio1_6_enable_vddio,
	input wire	gpio1_6_vtrip_sel,
	input wire	[1:0]	gpio1_6_ib_mode_sel,
	input wire	gpio1_6_out,
	input wire	[1:0]	gpio1_6_slew_ctl,
	input wire	gpio1_6_analog_pol,
	input wire	gpio1_6_analog_sel,
	input wire	gpio1_6_hys_trim,
	input wire	gpio1_6_hld_ovr,
	output wire	gpio1_6_in_h,
	input wire	gpio1_6_enable_h,
	output wire	gpio1_6_in,
	input wire	gpio1_6_hld_h_n,
	input wire	gpio1_6_enable_vdda_h,
	input wire	gpio1_6_analog_en,
	input wire	gpio1_6_enable_inp_h,
	input wire	gpio1_6_enable_vswitch_h,
	inout wire	gpio1_6_pad_a_noesd_h,
	inout wire	gpio1_6_pad_a_esd_0_h,
	inout wire	gpio1_6_pad_a_esd_1_h,
	output wire	gpio1_6_zero,
	output wire	gpio1_6_one,
	output wire	gpio1_7_tie_hi_esd,
	input wire	[2:0]	gpio1_7_dm,
	input wire	gpio1_7_slow,
	input wire	gpio1_7_oe_n,
	output wire	gpio1_7_tie_lo_esd,
	input wire	gpio1_7_inp_dis,
	input wire	gpio1_7_enable_vddio,
	input wire	gpio1_7_vtrip_sel,
	input wire	[1:0]	gpio1_7_ib_mode_sel,
	input wire	gpio1_7_out,
	input wire	[1:0]	gpio1_7_slew_ctl,
	input wire	gpio1_7_analog_pol,
	input wire	gpio1_7_analog_sel,
	input wire	gpio1_7_hys_trim,
	input wire	gpio1_7_hld_ovr,
	output wire	gpio1_7_in_h,
	input wire	gpio1_7_enable_h,
	output wire	gpio1_7_in,
	input wire	gpio1_7_hld_h_n,
	input wire	gpio1_7_enable_vdda_h,
	input wire	gpio1_7_analog_en,
	input wire	gpio1_7_enable_inp_h,
	input wire	gpio1_7_enable_vswitch_h,
	inout wire	gpio1_7_pad_a_noesd_h,
	inout wire	gpio1_7_pad_a_esd_0_h,
	inout wire	gpio1_7_pad_a_esd_1_h,
	output wire	gpio1_7_zero,
	output wire	gpio1_7_one,
	output wire	gpio2_0_tie_lo_esd,
	output wire	gpio2_0_in,
	output wire	gpio2_0_tie_hi_esd,
	input wire	gpio2_0_enable_vddio,
	input wire	gpio2_0_slow,
	inout wire	gpio2_0_pad_a_esd_0_h,
	inout wire	gpio2_0_pad_a_esd_1_h,
	inout wire	gpio2_0_pad_a_noesd_h,
	input wire	gpio2_0_analog_en,
	input wire	gpio2_0_analog_pol,
	input wire	gpio2_0_inp_dis,
	input wire	gpio2_0_enable_inp_h,
	input wire	gpio2_0_enable_h,
	input wire	gpio2_0_hld_h_n,
	input wire	gpio2_0_analog_sel,
	input wire	[2:0]	gpio2_0_dm,
	input wire	gpio2_0_hld_ovr,
	input wire	gpio2_0_out,
	input wire	gpio2_0_enable_vswitch_h,
	input wire	gpio2_0_enable_vdda_h,
	input wire	gpio2_0_vtrip_sel,
	input wire	gpio2_0_ib_mode_sel,
	input wire	gpio2_0_oe_n,
	output wire	gpio2_0_in_h,
	output wire	gpio2_0_zero,
	output wire	gpio2_0_one,
	output wire	gpio2_1_tie_lo_esd,
	output wire	gpio2_1_in,
	output wire	gpio2_1_tie_hi_esd,
	input wire	gpio2_1_enable_vddio,
	input wire	gpio2_1_slow,
	inout wire	gpio2_1_pad_a_esd_0_h,
	inout wire	gpio2_1_pad_a_esd_1_h,
	inout wire	gpio2_1_pad_a_noesd_h,
	input wire	gpio2_1_analog_en,
	input wire	gpio2_1_analog_pol,
	input wire	gpio2_1_inp_dis,
	input wire	gpio2_1_enable_inp_h,
	input wire	gpio2_1_enable_h,
	input wire	gpio2_1_hld_h_n,
	input wire	gpio2_1_analog_sel,
	input wire	[2:0]	gpio2_1_dm,
	input wire	gpio2_1_hld_ovr,
	input wire	gpio2_1_out,
	input wire	gpio2_1_enable_vswitch_h,
	input wire	gpio2_1_enable_vdda_h,
	input wire	gpio2_1_vtrip_sel,
	input wire	gpio2_1_ib_mode_sel,
	input wire	gpio2_1_oe_n,
	output wire	gpio2_1_in_h,
	output wire	gpio2_1_zero,
	output wire	gpio2_1_one,
	output wire	gpio2_2_tie_lo_esd,
	output wire	gpio2_2_in,
	output wire	gpio2_2_tie_hi_esd,
	input wire	gpio2_2_enable_vddio,
	input wire	gpio2_2_slow,
	inout wire	gpio2_2_pad_a_esd_0_h,
	inout wire	gpio2_2_pad_a_esd_1_h,
	inout wire	gpio2_2_pad_a_noesd_h,
	input wire	gpio2_2_analog_en,
	input wire	gpio2_2_analog_pol,
	input wire	gpio2_2_inp_dis,
	input wire	gpio2_2_enable_inp_h,
	input wire	gpio2_2_enable_h,
	input wire	gpio2_2_hld_h_n,
	input wire	gpio2_2_analog_sel,
	input wire	[2:0]	gpio2_2_dm,
	input wire	gpio2_2_hld_ovr,
	input wire	gpio2_2_out,
	input wire	gpio2_2_enable_vswitch_h,
	input wire	gpio2_2_enable_vdda_h,
	input wire	gpio2_2_vtrip_sel,
	input wire	gpio2_2_ib_mode_sel,
	input wire	gpio2_2_oe_n,
	output wire	gpio2_2_in_h,
	output wire	gpio2_2_zero,
	output wire	gpio2_2_one,
	output wire	gpio2_3_tie_lo_esd,
	output wire	gpio2_3_in,
	output wire	gpio2_3_tie_hi_esd,
	input wire	gpio2_3_enable_vddio,
	input wire	gpio2_3_slow,
	inout wire	gpio2_3_pad_a_esd_0_h,
	inout wire	gpio2_3_pad_a_esd_1_h,
	inout wire	gpio2_3_pad_a_noesd_h,
	input wire	gpio2_3_analog_en,
	input wire	gpio2_3_analog_pol,
	input wire	gpio2_3_inp_dis,
	input wire	gpio2_3_enable_inp_h,
	input wire	gpio2_3_enable_h,
	input wire	gpio2_3_hld_h_n,
	input wire	gpio2_3_analog_sel,
	input wire	[2:0]	gpio2_3_dm,
	input wire	gpio2_3_hld_ovr,
	input wire	gpio2_3_out,
	input wire	gpio2_3_enable_vswitch_h,
	input wire	gpio2_3_enable_vdda_h,
	input wire	gpio2_3_vtrip_sel,
	input wire	gpio2_3_ib_mode_sel,
	input wire	gpio2_3_oe_n,
	output wire	gpio2_3_in_h,
	output wire	gpio2_3_zero,
	output wire	gpio2_3_one,
	output wire	gpio2_4_tie_lo_esd,
	output wire	gpio2_4_in,
	output wire	gpio2_4_tie_hi_esd,
	input wire	gpio2_4_enable_vddio,
	input wire	gpio2_4_slow,
	inout wire	gpio2_4_pad_a_esd_0_h,
	inout wire	gpio2_4_pad_a_esd_1_h,
	inout wire	gpio2_4_pad_a_noesd_h,
	input wire	gpio2_4_analog_en,
	input wire	gpio2_4_analog_pol,
	input wire	gpio2_4_inp_dis,
	input wire	gpio2_4_enable_inp_h,
	input wire	gpio2_4_enable_h,
	input wire	gpio2_4_hld_h_n,
	input wire	gpio2_4_analog_sel,
	input wire	[2:0]	gpio2_4_dm,
	input wire	gpio2_4_hld_ovr,
	input wire	gpio2_4_out,
	input wire	gpio2_4_enable_vswitch_h,
	input wire	gpio2_4_enable_vdda_h,
	input wire	gpio2_4_vtrip_sel,
	input wire	gpio2_4_ib_mode_sel,
	input wire	gpio2_4_oe_n,
	output wire	gpio2_4_in_h,
	output wire	gpio2_4_zero,
	output wire	gpio2_4_one,
	output wire	gpio2_5_tie_lo_esd,
	output wire	gpio2_5_in,
	output wire	gpio2_5_tie_hi_esd,
	input wire	gpio2_5_enable_vddio,
	input wire	gpio2_5_slow,
	inout wire	gpio2_5_pad_a_esd_0_h,
	inout wire	gpio2_5_pad_a_esd_1_h,
	inout wire	gpio2_5_pad_a_noesd_h,
	input wire	gpio2_5_analog_en,
	input wire	gpio2_5_analog_pol,
	input wire	gpio2_5_inp_dis,
	input wire	gpio2_5_enable_inp_h,
	input wire	gpio2_5_enable_h,
	input wire	gpio2_5_hld_h_n,
	input wire	gpio2_5_analog_sel,
	input wire	[2:0]	gpio2_5_dm,
	input wire	gpio2_5_hld_ovr,
	input wire	gpio2_5_out,
	input wire	gpio2_5_enable_vswitch_h,
	input wire	gpio2_5_enable_vdda_h,
	input wire	gpio2_5_vtrip_sel,
	input wire	gpio2_5_ib_mode_sel,
	input wire	gpio2_5_oe_n,
	output wire	gpio2_5_in_h,
	output wire	gpio2_5_zero,
	output wire	gpio2_5_one,
	output wire	gpio2_6_tie_lo_esd,
	output wire	gpio2_6_in,
	output wire	gpio2_6_tie_hi_esd,
	input wire	gpio2_6_enable_vddio,
	input wire	gpio2_6_slow,
	inout wire	gpio2_6_pad_a_esd_0_h,
	inout wire	gpio2_6_pad_a_esd_1_h,
	inout wire	gpio2_6_pad_a_noesd_h,
	input wire	gpio2_6_analog_en,
	input wire	gpio2_6_analog_pol,
	input wire	gpio2_6_inp_dis,
	input wire	gpio2_6_enable_inp_h,
	input wire	gpio2_6_enable_h,
	input wire	gpio2_6_hld_h_n,
	input wire	gpio2_6_analog_sel,
	input wire	[2:0]	gpio2_6_dm,
	input wire	gpio2_6_hld_ovr,
	input wire	gpio2_6_out,
	input wire	gpio2_6_enable_vswitch_h,
	input wire	gpio2_6_enable_vdda_h,
	input wire	gpio2_6_vtrip_sel,
	input wire	gpio2_6_ib_mode_sel,
	input wire	gpio2_6_oe_n,
	output wire	gpio2_6_in_h,
	output wire	gpio2_6_zero,
	output wire	gpio2_6_one,
	output wire	gpio2_7_tie_lo_esd,
	output wire	gpio2_7_in,
	output wire	gpio2_7_tie_hi_esd,
	input wire	gpio2_7_enable_vddio,
	input wire	gpio2_7_slow,
	inout wire	gpio2_7_pad_a_esd_0_h,
	inout wire	gpio2_7_pad_a_esd_1_h,
	inout wire	gpio2_7_pad_a_noesd_h,
	input wire	gpio2_7_analog_en,
	input wire	gpio2_7_analog_pol,
	input wire	gpio2_7_inp_dis,
	input wire	gpio2_7_enable_inp_h,
	input wire	gpio2_7_enable_h,
	input wire	gpio2_7_hld_h_n,
	input wire	gpio2_7_analog_sel,
	input wire	[2:0]	gpio2_7_dm,
	input wire	gpio2_7_hld_ovr,
	input wire	gpio2_7_out,
	input wire	gpio2_7_enable_vswitch_h,
	input wire	gpio2_7_enable_vdda_h,
	input wire	gpio2_7_vtrip_sel,
	input wire	gpio2_7_ib_mode_sel,
	input wire	gpio2_7_oe_n,
	output wire	gpio2_7_in_h,
	output wire	gpio2_7_zero,
	output wire	gpio2_7_one,
	input wire	muxsplit_ne_hld_vdda_h_n,
	input wire	muxsplit_ne_enable_vdda_h,
	input wire	muxsplit_ne_switch_aa_sl,
	input wire	muxsplit_ne_switch_aa_s0,
	input wire	muxsplit_ne_switch_bb_s0,
	input wire	muxsplit_ne_switch_bb_sl,
	input wire	muxsplit_ne_switch_bb_sr,
	input wire	muxsplit_ne_switch_aa_sr,
	output wire	gpio3_0_tie_lo_esd,
	output wire	gpio3_0_in,
	output wire	gpio3_0_tie_hi_esd,
	input wire	gpio3_0_enable_vddio,
	input wire	gpio3_0_slow,
	inout wire	gpio3_0_pad_a_esd_0_h,
	inout wire	gpio3_0_pad_a_esd_1_h,
	inout wire	gpio3_0_pad_a_noesd_h,
	input wire	gpio3_0_analog_en,
	input wire	gpio3_0_analog_pol,
	input wire	gpio3_0_inp_dis,
	input wire	gpio3_0_enable_inp_h,
	input wire	gpio3_0_enable_h,
	input wire	gpio3_0_hld_h_n,
	input wire	gpio3_0_analog_sel,
	input wire	[2:0]	gpio3_0_dm,
	input wire	gpio3_0_hld_ovr,
	input wire	gpio3_0_out,
	input wire	gpio3_0_enable_vswitch_h,
	input wire	gpio3_0_enable_vdda_h,
	input wire	gpio3_0_vtrip_sel,
	input wire	gpio3_0_ib_mode_sel,
	input wire	gpio3_0_oe_n,
	output wire	gpio3_0_in_h,
	output wire	gpio3_0_zero,
	output wire	gpio3_0_one,
	output wire	gpio3_1_tie_lo_esd,
	output wire	gpio3_1_in,
	output wire	gpio3_1_tie_hi_esd,
	input wire	gpio3_1_enable_vddio,
	input wire	gpio3_1_slow,
	inout wire	gpio3_1_pad_a_esd_0_h,
	inout wire	gpio3_1_pad_a_esd_1_h,
	inout wire	gpio3_1_pad_a_noesd_h,
	input wire	gpio3_1_analog_en,
	input wire	gpio3_1_analog_pol,
	input wire	gpio3_1_inp_dis,
	input wire	gpio3_1_enable_inp_h,
	input wire	gpio3_1_enable_h,
	input wire	gpio3_1_hld_h_n,
	input wire	gpio3_1_analog_sel,
	input wire	[2:0]	gpio3_1_dm,
	input wire	gpio3_1_hld_ovr,
	input wire	gpio3_1_out,
	input wire	gpio3_1_enable_vswitch_h,
	input wire	gpio3_1_enable_vdda_h,
	input wire	gpio3_1_vtrip_sel,
	input wire	gpio3_1_ib_mode_sel,
	input wire	gpio3_1_oe_n,
	output wire	gpio3_1_in_h,
	output wire	gpio3_1_zero,
	output wire	gpio3_1_one,
	output wire	gpio3_2_tie_lo_esd,
	output wire	gpio3_2_in,
	output wire	gpio3_2_tie_hi_esd,
	input wire	gpio3_2_enable_vddio,
	input wire	gpio3_2_slow,
	inout wire	gpio3_2_pad_a_esd_0_h,
	inout wire	gpio3_2_pad_a_esd_1_h,
	inout wire	gpio3_2_pad_a_noesd_h,
	input wire	gpio3_2_analog_en,
	input wire	gpio3_2_analog_pol,
	input wire	gpio3_2_inp_dis,
	input wire	gpio3_2_enable_inp_h,
	input wire	gpio3_2_enable_h,
	input wire	gpio3_2_hld_h_n,
	input wire	gpio3_2_analog_sel,
	input wire	[2:0]	gpio3_2_dm,
	input wire	gpio3_2_hld_ovr,
	input wire	gpio3_2_out,
	input wire	gpio3_2_enable_vswitch_h,
	input wire	gpio3_2_enable_vdda_h,
	input wire	gpio3_2_vtrip_sel,
	input wire	gpio3_2_ib_mode_sel,
	input wire	gpio3_2_oe_n,
	output wire	gpio3_2_in_h,
	output wire	gpio3_2_zero,
	output wire	gpio3_2_one,
	output wire	gpio3_3_tie_lo_esd,
	output wire	gpio3_3_in,
	output wire	gpio3_3_tie_hi_esd,
	input wire	gpio3_3_enable_vddio,
	input wire	gpio3_3_slow,
	inout wire	gpio3_3_pad_a_esd_0_h,
	inout wire	gpio3_3_pad_a_esd_1_h,
	inout wire	gpio3_3_pad_a_noesd_h,
	input wire	gpio3_3_analog_en,
	input wire	gpio3_3_analog_pol,
	input wire	gpio3_3_inp_dis,
	input wire	gpio3_3_enable_inp_h,
	input wire	gpio3_3_enable_h,
	input wire	gpio3_3_hld_h_n,
	input wire	gpio3_3_analog_sel,
	input wire	[2:0]	gpio3_3_dm,
	input wire	gpio3_3_hld_ovr,
	input wire	gpio3_3_out,
	input wire	gpio3_3_enable_vswitch_h,
	input wire	gpio3_3_enable_vdda_h,
	input wire	gpio3_3_vtrip_sel,
	input wire	gpio3_3_ib_mode_sel,
	input wire	gpio3_3_oe_n,
	output wire	gpio3_3_in_h,
	output wire	gpio3_3_zero,
	output wire	gpio3_3_one,
	output wire	gpio3_4_tie_lo_esd,
	output wire	gpio3_4_in,
	output wire	gpio3_4_tie_hi_esd,
	input wire	gpio3_4_enable_vddio,
	input wire	gpio3_4_slow,
	inout wire	gpio3_4_pad_a_esd_0_h,
	inout wire	gpio3_4_pad_a_esd_1_h,
	inout wire	gpio3_4_pad_a_noesd_h,
	input wire	gpio3_4_analog_en,
	input wire	gpio3_4_analog_pol,
	input wire	gpio3_4_inp_dis,
	input wire	gpio3_4_enable_inp_h,
	input wire	gpio3_4_enable_h,
	input wire	gpio3_4_hld_h_n,
	input wire	gpio3_4_analog_sel,
	input wire	[2:0]	gpio3_4_dm,
	input wire	gpio3_4_hld_ovr,
	input wire	gpio3_4_out,
	input wire	gpio3_4_enable_vswitch_h,
	input wire	gpio3_4_enable_vdda_h,
	input wire	gpio3_4_vtrip_sel,
	input wire	gpio3_4_ib_mode_sel,
	input wire	gpio3_4_oe_n,
	output wire	gpio3_4_in_h,
	output wire	gpio3_4_zero,
	output wire	gpio3_4_one,
	output wire	gpio3_5_tie_lo_esd,
	output wire	gpio3_5_in,
	output wire	gpio3_5_tie_hi_esd,
	input wire	gpio3_5_enable_vddio,
	input wire	gpio3_5_slow,
	inout wire	gpio3_5_pad_a_esd_0_h,
	inout wire	gpio3_5_pad_a_esd_1_h,
	inout wire	gpio3_5_pad_a_noesd_h,
	input wire	gpio3_5_analog_en,
	input wire	gpio3_5_analog_pol,
	input wire	gpio3_5_inp_dis,
	input wire	gpio3_5_enable_inp_h,
	input wire	gpio3_5_enable_h,
	input wire	gpio3_5_hld_h_n,
	input wire	gpio3_5_analog_sel,
	input wire	[2:0]	gpio3_5_dm,
	input wire	gpio3_5_hld_ovr,
	input wire	gpio3_5_out,
	input wire	gpio3_5_enable_vswitch_h,
	input wire	gpio3_5_enable_vdda_h,
	input wire	gpio3_5_vtrip_sel,
	input wire	gpio3_5_ib_mode_sel,
	input wire	gpio3_5_oe_n,
	output wire	gpio3_5_in_h,
	output wire	gpio3_5_zero,
	output wire	gpio3_5_one,
	output wire	gpio3_6_tie_lo_esd,
	output wire	gpio3_6_in,
	output wire	gpio3_6_tie_hi_esd,
	input wire	gpio3_6_enable_vddio,
	input wire	gpio3_6_slow,
	inout wire	gpio3_6_pad_a_esd_0_h,
	inout wire	gpio3_6_pad_a_esd_1_h,
	inout wire	gpio3_6_pad_a_noesd_h,
	input wire	gpio3_6_analog_en,
	input wire	gpio3_6_analog_pol,
	input wire	gpio3_6_inp_dis,
	input wire	gpio3_6_enable_inp_h,
	input wire	gpio3_6_enable_h,
	input wire	gpio3_6_hld_h_n,
	input wire	gpio3_6_analog_sel,
	input wire	[2:0]	gpio3_6_dm,
	input wire	gpio3_6_hld_ovr,
	input wire	gpio3_6_out,
	input wire	gpio3_6_enable_vswitch_h,
	input wire	gpio3_6_enable_vdda_h,
	input wire	gpio3_6_vtrip_sel,
	input wire	gpio3_6_ib_mode_sel,
	input wire	gpio3_6_oe_n,
	output wire	gpio3_6_in_h,
	output wire	gpio3_6_zero,
	output wire	gpio3_6_one,
	output wire	gpio3_7_tie_lo_esd,
	output wire	gpio3_7_in,
	output wire	gpio3_7_tie_hi_esd,
	input wire	gpio3_7_enable_vddio,
	input wire	gpio3_7_slow,
	inout wire	gpio3_7_pad_a_esd_0_h,
	inout wire	gpio3_7_pad_a_esd_1_h,
	inout wire	gpio3_7_pad_a_noesd_h,
	input wire	gpio3_7_analog_en,
	input wire	gpio3_7_analog_pol,
	input wire	gpio3_7_inp_dis,
	input wire	gpio3_7_enable_inp_h,
	input wire	gpio3_7_enable_h,
	input wire	gpio3_7_hld_h_n,
	input wire	gpio3_7_analog_sel,
	input wire	[2:0]	gpio3_7_dm,
	input wire	gpio3_7_hld_ovr,
	input wire	gpio3_7_out,
	input wire	gpio3_7_enable_vswitch_h,
	input wire	gpio3_7_enable_vdda_h,
	input wire	gpio3_7_vtrip_sel,
	input wire	gpio3_7_ib_mode_sel,
	input wire	gpio3_7_oe_n,
	output wire	gpio3_7_in_h,
	output wire	gpio3_7_zero,
	output wire	gpio3_7_one,
	inout wire	analog_0_core,
	inout wire	analog_1_core,
	output wire	gpio4_0_tie_lo_esd,
	output wire	gpio4_0_in,
	output wire	gpio4_0_tie_hi_esd,
	input wire	gpio4_0_enable_vddio,
	input wire	gpio4_0_slow,
	inout wire	gpio4_0_pad_a_esd_0_h,
	inout wire	gpio4_0_pad_a_esd_1_h,
	inout wire	gpio4_0_pad_a_noesd_h,
	input wire	gpio4_0_analog_en,
	input wire	gpio4_0_analog_pol,
	input wire	gpio4_0_inp_dis,
	input wire	gpio4_0_enable_inp_h,
	input wire	gpio4_0_enable_h,
	input wire	gpio4_0_hld_h_n,
	input wire	gpio4_0_analog_sel,
	input wire	[2:0]	gpio4_0_dm,
	input wire	gpio4_0_hld_ovr,
	input wire	gpio4_0_out,
	input wire	gpio4_0_enable_vswitch_h,
	input wire	gpio4_0_enable_vdda_h,
	input wire	gpio4_0_vtrip_sel,
	input wire	gpio4_0_ib_mode_sel,
	input wire	gpio4_0_oe_n,
	output wire	gpio4_0_in_h,
	output wire	gpio4_0_zero,
	output wire	gpio4_0_one,
	output wire	gpio4_1_tie_lo_esd,
	output wire	gpio4_1_in,
	output wire	gpio4_1_tie_hi_esd,
	input wire	gpio4_1_enable_vddio,
	input wire	gpio4_1_slow,
	inout wire	gpio4_1_pad_a_esd_0_h,
	inout wire	gpio4_1_pad_a_esd_1_h,
	inout wire	gpio4_1_pad_a_noesd_h,
	input wire	gpio4_1_analog_en,
	input wire	gpio4_1_analog_pol,
	input wire	gpio4_1_inp_dis,
	input wire	gpio4_1_enable_inp_h,
	input wire	gpio4_1_enable_h,
	input wire	gpio4_1_hld_h_n,
	input wire	gpio4_1_analog_sel,
	input wire	[2:0]	gpio4_1_dm,
	input wire	gpio4_1_hld_ovr,
	input wire	gpio4_1_out,
	input wire	gpio4_1_enable_vswitch_h,
	input wire	gpio4_1_enable_vdda_h,
	input wire	gpio4_1_vtrip_sel,
	input wire	gpio4_1_ib_mode_sel,
	input wire	gpio4_1_oe_n,
	output wire	gpio4_1_in_h,
	output wire	gpio4_1_zero,
	output wire	gpio4_1_one,
	output wire	gpio4_2_tie_lo_esd,
	output wire	gpio4_2_in,
	output wire	gpio4_2_tie_hi_esd,
	input wire	gpio4_2_enable_vddio,
	input wire	gpio4_2_slow,
	inout wire	gpio4_2_pad_a_esd_0_h,
	inout wire	gpio4_2_pad_a_esd_1_h,
	inout wire	gpio4_2_pad_a_noesd_h,
	input wire	gpio4_2_analog_en,
	input wire	gpio4_2_analog_pol,
	input wire	gpio4_2_inp_dis,
	input wire	gpio4_2_enable_inp_h,
	input wire	gpio4_2_enable_h,
	input wire	gpio4_2_hld_h_n,
	input wire	gpio4_2_analog_sel,
	input wire	[2:0]	gpio4_2_dm,
	input wire	gpio4_2_hld_ovr,
	input wire	gpio4_2_out,
	input wire	gpio4_2_enable_vswitch_h,
	input wire	gpio4_2_enable_vdda_h,
	input wire	gpio4_2_vtrip_sel,
	input wire	gpio4_2_ib_mode_sel,
	input wire	gpio4_2_oe_n,
	output wire	gpio4_2_in_h,
	output wire	gpio4_2_zero,
	output wire	gpio4_2_one,
	output wire	gpio4_3_tie_lo_esd,
	output wire	gpio4_3_in,
	output wire	gpio4_3_tie_hi_esd,
	input wire	gpio4_3_enable_vddio,
	input wire	gpio4_3_slow,
	inout wire	gpio4_3_pad_a_esd_0_h,
	inout wire	gpio4_3_pad_a_esd_1_h,
	inout wire	gpio4_3_pad_a_noesd_h,
	input wire	gpio4_3_analog_en,
	input wire	gpio4_3_analog_pol,
	input wire	gpio4_3_inp_dis,
	input wire	gpio4_3_enable_inp_h,
	input wire	gpio4_3_enable_h,
	input wire	gpio4_3_hld_h_n,
	input wire	gpio4_3_analog_sel,
	input wire	[2:0]	gpio4_3_dm,
	input wire	gpio4_3_hld_ovr,
	input wire	gpio4_3_out,
	input wire	gpio4_3_enable_vswitch_h,
	input wire	gpio4_3_enable_vdda_h,
	input wire	gpio4_3_vtrip_sel,
	input wire	gpio4_3_ib_mode_sel,
	input wire	gpio4_3_oe_n,
	output wire	gpio4_3_in_h,
	output wire	gpio4_3_zero,
	output wire	gpio4_3_one,
	output wire	gpio4_4_tie_lo_esd,
	output wire	gpio4_4_in,
	output wire	gpio4_4_tie_hi_esd,
	input wire	gpio4_4_enable_vddio,
	input wire	gpio4_4_slow,
	inout wire	gpio4_4_pad_a_esd_0_h,
	inout wire	gpio4_4_pad_a_esd_1_h,
	inout wire	gpio4_4_pad_a_noesd_h,
	input wire	gpio4_4_analog_en,
	input wire	gpio4_4_analog_pol,
	input wire	gpio4_4_inp_dis,
	input wire	gpio4_4_enable_inp_h,
	input wire	gpio4_4_enable_h,
	input wire	gpio4_4_hld_h_n,
	input wire	gpio4_4_analog_sel,
	input wire	[2:0]	gpio4_4_dm,
	input wire	gpio4_4_hld_ovr,
	input wire	gpio4_4_out,
	input wire	gpio4_4_enable_vswitch_h,
	input wire	gpio4_4_enable_vdda_h,
	input wire	gpio4_4_vtrip_sel,
	input wire	gpio4_4_ib_mode_sel,
	input wire	gpio4_4_oe_n,
	output wire	gpio4_4_in_h,
	output wire	gpio4_4_zero,
	output wire	gpio4_4_one,
	output wire	gpio4_5_tie_lo_esd,
	output wire	gpio4_5_in,
	output wire	gpio4_5_tie_hi_esd,
	input wire	gpio4_5_enable_vddio,
	input wire	gpio4_5_slow,
	inout wire	gpio4_5_pad_a_esd_0_h,
	inout wire	gpio4_5_pad_a_esd_1_h,
	inout wire	gpio4_5_pad_a_noesd_h,
	input wire	gpio4_5_analog_en,
	input wire	gpio4_5_analog_pol,
	input wire	gpio4_5_inp_dis,
	input wire	gpio4_5_enable_inp_h,
	input wire	gpio4_5_enable_h,
	input wire	gpio4_5_hld_h_n,
	input wire	gpio4_5_analog_sel,
	input wire	[2:0]	gpio4_5_dm,
	input wire	gpio4_5_hld_ovr,
	input wire	gpio4_5_out,
	input wire	gpio4_5_enable_vswitch_h,
	input wire	gpio4_5_enable_vdda_h,
	input wire	gpio4_5_vtrip_sel,
	input wire	gpio4_5_ib_mode_sel,
	input wire	gpio4_5_oe_n,
	output wire	gpio4_5_in_h,
	output wire	gpio4_5_zero,
	output wire	gpio4_5_one,
	output wire	gpio4_6_tie_lo_esd,
	output wire	gpio4_6_in,
	output wire	gpio4_6_tie_hi_esd,
	input wire	gpio4_6_enable_vddio,
	input wire	gpio4_6_slow,
	inout wire	gpio4_6_pad_a_esd_0_h,
	inout wire	gpio4_6_pad_a_esd_1_h,
	inout wire	gpio4_6_pad_a_noesd_h,
	input wire	gpio4_6_analog_en,
	input wire	gpio4_6_analog_pol,
	input wire	gpio4_6_inp_dis,
	input wire	gpio4_6_enable_inp_h,
	input wire	gpio4_6_enable_h,
	input wire	gpio4_6_hld_h_n,
	input wire	gpio4_6_analog_sel,
	input wire	[2:0]	gpio4_6_dm,
	input wire	gpio4_6_hld_ovr,
	input wire	gpio4_6_out,
	input wire	gpio4_6_enable_vswitch_h,
	input wire	gpio4_6_enable_vdda_h,
	input wire	gpio4_6_vtrip_sel,
	input wire	gpio4_6_ib_mode_sel,
	input wire	gpio4_6_oe_n,
	output wire	gpio4_6_in_h,
	output wire	gpio4_6_zero,
	output wire	gpio4_6_one,
	output wire	gpio4_7_tie_lo_esd,
	output wire	gpio4_7_in,
	output wire	gpio4_7_tie_hi_esd,
	input wire	gpio4_7_enable_vddio,
	input wire	gpio4_7_slow,
	inout wire	gpio4_7_pad_a_esd_0_h,
	inout wire	gpio4_7_pad_a_esd_1_h,
	inout wire	gpio4_7_pad_a_noesd_h,
	input wire	gpio4_7_analog_en,
	input wire	gpio4_7_analog_pol,
	input wire	gpio4_7_inp_dis,
	input wire	gpio4_7_enable_inp_h,
	input wire	gpio4_7_enable_h,
	input wire	gpio4_7_hld_h_n,
	input wire	gpio4_7_analog_sel,
	input wire	[2:0]	gpio4_7_dm,
	input wire	gpio4_7_hld_ovr,
	input wire	gpio4_7_out,
	input wire	gpio4_7_enable_vswitch_h,
	input wire	gpio4_7_enable_vdda_h,
	input wire	gpio4_7_vtrip_sel,
	input wire	gpio4_7_ib_mode_sel,
	input wire	gpio4_7_oe_n,
	output wire	gpio4_7_in_h,
	output wire	gpio4_7_zero,
	output wire	gpio4_7_one,
	input wire	muxsplit_nw_hld_vdda_h_n,
	input wire	muxsplit_nw_enable_vdda_h,
	input wire	muxsplit_nw_switch_aa_sl,
	input wire	muxsplit_nw_switch_aa_s0,
	input wire	muxsplit_nw_switch_bb_s0,
	input wire	muxsplit_nw_switch_bb_sl,
	input wire	muxsplit_nw_switch_bb_sr,
	input wire	muxsplit_nw_switch_aa_sr,
	output wire	gpio5_0_tie_lo_esd,
	output wire	gpio5_0_in,
	output wire	gpio5_0_tie_hi_esd,
	input wire	gpio5_0_enable_vddio,
	input wire	gpio5_0_slow,
	inout wire	gpio5_0_pad_a_esd_0_h,
	inout wire	gpio5_0_pad_a_esd_1_h,
	inout wire	gpio5_0_pad_a_noesd_h,
	input wire	gpio5_0_analog_en,
	input wire	gpio5_0_analog_pol,
	input wire	gpio5_0_inp_dis,
	input wire	gpio5_0_enable_inp_h,
	input wire	gpio5_0_enable_h,
	input wire	gpio5_0_hld_h_n,
	input wire	gpio5_0_analog_sel,
	input wire	[2:0]	gpio5_0_dm,
	input wire	gpio5_0_hld_ovr,
	input wire	gpio5_0_out,
	input wire	gpio5_0_enable_vswitch_h,
	input wire	gpio5_0_enable_vdda_h,
	input wire	gpio5_0_vtrip_sel,
	input wire	gpio5_0_ib_mode_sel,
	input wire	gpio5_0_oe_n,
	output wire	gpio5_0_in_h,
	output wire	gpio5_0_zero,
	output wire	gpio5_0_one,
	output wire	gpio5_1_tie_lo_esd,
	output wire	gpio5_1_in,
	output wire	gpio5_1_tie_hi_esd,
	input wire	gpio5_1_enable_vddio,
	input wire	gpio5_1_slow,
	inout wire	gpio5_1_pad_a_esd_0_h,
	inout wire	gpio5_1_pad_a_esd_1_h,
	inout wire	gpio5_1_pad_a_noesd_h,
	input wire	gpio5_1_analog_en,
	input wire	gpio5_1_analog_pol,
	input wire	gpio5_1_inp_dis,
	input wire	gpio5_1_enable_inp_h,
	input wire	gpio5_1_enable_h,
	input wire	gpio5_1_hld_h_n,
	input wire	gpio5_1_analog_sel,
	input wire	[2:0]	gpio5_1_dm,
	input wire	gpio5_1_hld_ovr,
	input wire	gpio5_1_out,
	input wire	gpio5_1_enable_vswitch_h,
	input wire	gpio5_1_enable_vdda_h,
	input wire	gpio5_1_vtrip_sel,
	input wire	gpio5_1_ib_mode_sel,
	input wire	gpio5_1_oe_n,
	output wire	gpio5_1_in_h,
	output wire	gpio5_1_zero,
	output wire	gpio5_1_one,
	output wire	gpio5_2_tie_lo_esd,
	output wire	gpio5_2_in,
	output wire	gpio5_2_tie_hi_esd,
	input wire	gpio5_2_enable_vddio,
	input wire	gpio5_2_slow,
	inout wire	gpio5_2_pad_a_esd_0_h,
	inout wire	gpio5_2_pad_a_esd_1_h,
	inout wire	gpio5_2_pad_a_noesd_h,
	input wire	gpio5_2_analog_en,
	input wire	gpio5_2_analog_pol,
	input wire	gpio5_2_inp_dis,
	input wire	gpio5_2_enable_inp_h,
	input wire	gpio5_2_enable_h,
	input wire	gpio5_2_hld_h_n,
	input wire	gpio5_2_analog_sel,
	input wire	[2:0]	gpio5_2_dm,
	input wire	gpio5_2_hld_ovr,
	input wire	gpio5_2_out,
	input wire	gpio5_2_enable_vswitch_h,
	input wire	gpio5_2_enable_vdda_h,
	input wire	gpio5_2_vtrip_sel,
	input wire	gpio5_2_ib_mode_sel,
	input wire	gpio5_2_oe_n,
	output wire	gpio5_2_in_h,
	output wire	gpio5_2_zero,
	output wire	gpio5_2_one,
	output wire	gpio5_3_tie_lo_esd,
	output wire	gpio5_3_in,
	output wire	gpio5_3_tie_hi_esd,
	input wire	gpio5_3_enable_vddio,
	input wire	gpio5_3_slow,
	inout wire	gpio5_3_pad_a_esd_0_h,
	inout wire	gpio5_3_pad_a_esd_1_h,
	inout wire	gpio5_3_pad_a_noesd_h,
	input wire	gpio5_3_analog_en,
	input wire	gpio5_3_analog_pol,
	input wire	gpio5_3_inp_dis,
	input wire	gpio5_3_enable_inp_h,
	input wire	gpio5_3_enable_h,
	input wire	gpio5_3_hld_h_n,
	input wire	gpio5_3_analog_sel,
	input wire	[2:0]	gpio5_3_dm,
	input wire	gpio5_3_hld_ovr,
	input wire	gpio5_3_out,
	input wire	gpio5_3_enable_vswitch_h,
	input wire	gpio5_3_enable_vdda_h,
	input wire	gpio5_3_vtrip_sel,
	input wire	gpio5_3_ib_mode_sel,
	input wire	gpio5_3_oe_n,
	output wire	gpio5_3_in_h,
	output wire	gpio5_3_zero,
	output wire	gpio5_3_one,
	output wire	gpio5_4_tie_lo_esd,
	output wire	gpio5_4_in,
	output wire	gpio5_4_tie_hi_esd,
	input wire	gpio5_4_enable_vddio,
	input wire	gpio5_4_slow,
	inout wire	gpio5_4_pad_a_esd_0_h,
	inout wire	gpio5_4_pad_a_esd_1_h,
	inout wire	gpio5_4_pad_a_noesd_h,
	input wire	gpio5_4_analog_en,
	input wire	gpio5_4_analog_pol,
	input wire	gpio5_4_inp_dis,
	input wire	gpio5_4_enable_inp_h,
	input wire	gpio5_4_enable_h,
	input wire	gpio5_4_hld_h_n,
	input wire	gpio5_4_analog_sel,
	input wire	[2:0]	gpio5_4_dm,
	input wire	gpio5_4_hld_ovr,
	input wire	gpio5_4_out,
	input wire	gpio5_4_enable_vswitch_h,
	input wire	gpio5_4_enable_vdda_h,
	input wire	gpio5_4_vtrip_sel,
	input wire	gpio5_4_ib_mode_sel,
	input wire	gpio5_4_oe_n,
	output wire	gpio5_4_in_h,
	output wire	gpio5_4_zero,
	output wire	gpio5_4_one,
	output wire	gpio5_5_tie_lo_esd,
	output wire	gpio5_5_in,
	output wire	gpio5_5_tie_hi_esd,
	input wire	gpio5_5_enable_vddio,
	input wire	gpio5_5_slow,
	inout wire	gpio5_5_pad_a_esd_0_h,
	inout wire	gpio5_5_pad_a_esd_1_h,
	inout wire	gpio5_5_pad_a_noesd_h,
	input wire	gpio5_5_analog_en,
	input wire	gpio5_5_analog_pol,
	input wire	gpio5_5_inp_dis,
	input wire	gpio5_5_enable_inp_h,
	input wire	gpio5_5_enable_h,
	input wire	gpio5_5_hld_h_n,
	input wire	gpio5_5_analog_sel,
	input wire	[2:0]	gpio5_5_dm,
	input wire	gpio5_5_hld_ovr,
	input wire	gpio5_5_out,
	input wire	gpio5_5_enable_vswitch_h,
	input wire	gpio5_5_enable_vdda_h,
	input wire	gpio5_5_vtrip_sel,
	input wire	gpio5_5_ib_mode_sel,
	input wire	gpio5_5_oe_n,
	output wire	gpio5_5_in_h,
	output wire	gpio5_5_zero,
	output wire	gpio5_5_one,
	output wire	gpio5_6_tie_lo_esd,
	output wire	gpio5_6_in,
	output wire	gpio5_6_tie_hi_esd,
	input wire	gpio5_6_enable_vddio,
	input wire	gpio5_6_slow,
	inout wire	gpio5_6_pad_a_esd_0_h,
	inout wire	gpio5_6_pad_a_esd_1_h,
	inout wire	gpio5_6_pad_a_noesd_h,
	input wire	gpio5_6_analog_en,
	input wire	gpio5_6_analog_pol,
	input wire	gpio5_6_inp_dis,
	input wire	gpio5_6_enable_inp_h,
	input wire	gpio5_6_enable_h,
	input wire	gpio5_6_hld_h_n,
	input wire	gpio5_6_analog_sel,
	input wire	[2:0]	gpio5_6_dm,
	input wire	gpio5_6_hld_ovr,
	input wire	gpio5_6_out,
	input wire	gpio5_6_enable_vswitch_h,
	input wire	gpio5_6_enable_vdda_h,
	input wire	gpio5_6_vtrip_sel,
	input wire	gpio5_6_ib_mode_sel,
	input wire	gpio5_6_oe_n,
	output wire	gpio5_6_in_h,
	output wire	gpio5_6_zero,
	output wire	gpio5_6_one,
	output wire	gpio5_7_tie_lo_esd,
	output wire	gpio5_7_in,
	output wire	gpio5_7_tie_hi_esd,
	input wire	gpio5_7_enable_vddio,
	input wire	gpio5_7_slow,
	inout wire	gpio5_7_pad_a_esd_0_h,
	inout wire	gpio5_7_pad_a_esd_1_h,
	inout wire	gpio5_7_pad_a_noesd_h,
	input wire	gpio5_7_analog_en,
	input wire	gpio5_7_analog_pol,
	input wire	gpio5_7_inp_dis,
	input wire	gpio5_7_enable_inp_h,
	input wire	gpio5_7_enable_h,
	input wire	gpio5_7_hld_h_n,
	input wire	gpio5_7_analog_sel,
	input wire	[2:0]	gpio5_7_dm,
	input wire	gpio5_7_hld_ovr,
	input wire	gpio5_7_out,
	input wire	gpio5_7_enable_vswitch_h,
	input wire	gpio5_7_enable_vdda_h,
	input wire	gpio5_7_vtrip_sel,
	input wire	gpio5_7_ib_mode_sel,
	input wire	gpio5_7_oe_n,
	output wire	gpio5_7_in_h,
	output wire	gpio5_7_zero,
	output wire	gpio5_7_one,
	output wire	gpio6_0_tie_hi_esd,
	input wire	[2:0]	gpio6_0_dm,
	input wire	gpio6_0_slow,
	input wire	gpio6_0_oe_n,
	output wire	gpio6_0_tie_lo_esd,
	input wire	gpio6_0_inp_dis,
	input wire	gpio6_0_enable_vddio,
	input wire	gpio6_0_vtrip_sel,
	input wire	[1:0]	gpio6_0_ib_mode_sel,
	input wire	gpio6_0_out,
	input wire	[1:0]	gpio6_0_slew_ctl,
	input wire	gpio6_0_analog_pol,
	input wire	gpio6_0_analog_sel,
	input wire	gpio6_0_hys_trim,
	input wire	gpio6_0_hld_ovr,
	output wire	gpio6_0_in_h,
	input wire	gpio6_0_enable_h,
	output wire	gpio6_0_in,
	input wire	gpio6_0_hld_h_n,
	input wire	gpio6_0_enable_vdda_h,
	input wire	gpio6_0_analog_en,
	input wire	gpio6_0_enable_inp_h,
	input wire	gpio6_0_enable_vswitch_h,
	inout wire	gpio6_0_pad_a_noesd_h,
	inout wire	gpio6_0_pad_a_esd_0_h,
	inout wire	gpio6_0_pad_a_esd_1_h,
	output wire	gpio6_0_zero,
	output wire	gpio6_0_one,
	output wire	gpio6_1_tie_hi_esd,
	input wire	[2:0]	gpio6_1_dm,
	input wire	gpio6_1_slow,
	input wire	gpio6_1_oe_n,
	output wire	gpio6_1_tie_lo_esd,
	input wire	gpio6_1_inp_dis,
	input wire	gpio6_1_enable_vddio,
	input wire	gpio6_1_vtrip_sel,
	input wire	[1:0]	gpio6_1_ib_mode_sel,
	input wire	gpio6_1_out,
	input wire	[1:0]	gpio6_1_slew_ctl,
	input wire	gpio6_1_analog_pol,
	input wire	gpio6_1_analog_sel,
	input wire	gpio6_1_hys_trim,
	input wire	gpio6_1_hld_ovr,
	output wire	gpio6_1_in_h,
	input wire	gpio6_1_enable_h,
	output wire	gpio6_1_in,
	input wire	gpio6_1_hld_h_n,
	input wire	gpio6_1_enable_vdda_h,
	input wire	gpio6_1_analog_en,
	input wire	gpio6_1_enable_inp_h,
	input wire	gpio6_1_enable_vswitch_h,
	inout wire	gpio6_1_pad_a_noesd_h,
	inout wire	gpio6_1_pad_a_esd_0_h,
	inout wire	gpio6_1_pad_a_esd_1_h,
	output wire	gpio6_1_zero,
	output wire	gpio6_1_one,
	output wire	gpio6_2_tie_hi_esd,
	input wire	[2:0]	gpio6_2_dm,
	input wire	gpio6_2_slow,
	input wire	gpio6_2_oe_n,
	output wire	gpio6_2_tie_lo_esd,
	input wire	gpio6_2_inp_dis,
	input wire	gpio6_2_enable_vddio,
	input wire	gpio6_2_vtrip_sel,
	input wire	[1:0]	gpio6_2_ib_mode_sel,
	input wire	gpio6_2_out,
	input wire	[1:0]	gpio6_2_slew_ctl,
	input wire	gpio6_2_analog_pol,
	input wire	gpio6_2_analog_sel,
	input wire	gpio6_2_hys_trim,
	input wire	gpio6_2_hld_ovr,
	output wire	gpio6_2_in_h,
	input wire	gpio6_2_enable_h,
	output wire	gpio6_2_in,
	input wire	gpio6_2_hld_h_n,
	input wire	gpio6_2_enable_vdda_h,
	input wire	gpio6_2_analog_en,
	input wire	gpio6_2_enable_inp_h,
	input wire	gpio6_2_enable_vswitch_h,
	inout wire	gpio6_2_pad_a_noesd_h,
	inout wire	gpio6_2_pad_a_esd_0_h,
	inout wire	gpio6_2_pad_a_esd_1_h,
	output wire	gpio6_2_zero,
	output wire	gpio6_2_one,
	output wire	gpio6_3_tie_hi_esd,
	input wire	[2:0]	gpio6_3_dm,
	input wire	gpio6_3_slow,
	input wire	gpio6_3_oe_n,
	output wire	gpio6_3_tie_lo_esd,
	input wire	gpio6_3_inp_dis,
	input wire	gpio6_3_enable_vddio,
	input wire	gpio6_3_vtrip_sel,
	input wire	[1:0]	gpio6_3_ib_mode_sel,
	input wire	gpio6_3_out,
	input wire	[1:0]	gpio6_3_slew_ctl,
	input wire	gpio6_3_analog_pol,
	input wire	gpio6_3_analog_sel,
	input wire	gpio6_3_hys_trim,
	input wire	gpio6_3_hld_ovr,
	output wire	gpio6_3_in_h,
	input wire	gpio6_3_enable_h,
	output wire	gpio6_3_in,
	input wire	gpio6_3_hld_h_n,
	input wire	gpio6_3_enable_vdda_h,
	input wire	gpio6_3_analog_en,
	input wire	gpio6_3_enable_inp_h,
	input wire	gpio6_3_enable_vswitch_h,
	inout wire	gpio6_3_pad_a_noesd_h,
	inout wire	gpio6_3_pad_a_esd_0_h,
	inout wire	gpio6_3_pad_a_esd_1_h,
	output wire	gpio6_3_zero,
	output wire	gpio6_3_one,
	input wire	[4:0]	vref_w_ref_sel,
	inout wire	vref_w_vinref,
	input wire	vref_w_enable_h,
	input wire	vref_w_hld_h_n,
	input wire	vref_w_vrefgen_en,
	output wire	gpio6_4_tie_hi_esd,
	input wire	[2:0]	gpio6_4_dm,
	input wire	gpio6_4_slow,
	input wire	gpio6_4_oe_n,
	output wire	gpio6_4_tie_lo_esd,
	input wire	gpio6_4_inp_dis,
	input wire	gpio6_4_enable_vddio,
	input wire	gpio6_4_vtrip_sel,
	input wire	[1:0]	gpio6_4_ib_mode_sel,
	input wire	gpio6_4_out,
	input wire	[1:0]	gpio6_4_slew_ctl,
	input wire	gpio6_4_analog_pol,
	input wire	gpio6_4_analog_sel,
	input wire	gpio6_4_hys_trim,
	input wire	gpio6_4_hld_ovr,
	output wire	gpio6_4_in_h,
	input wire	gpio6_4_enable_h,
	output wire	gpio6_4_in,
	input wire	gpio6_4_hld_h_n,
	input wire	gpio6_4_enable_vdda_h,
	input wire	gpio6_4_analog_en,
	input wire	gpio6_4_enable_inp_h,
	input wire	gpio6_4_enable_vswitch_h,
	inout wire	gpio6_4_pad_a_noesd_h,
	inout wire	gpio6_4_pad_a_esd_0_h,
	inout wire	gpio6_4_pad_a_esd_1_h,
	output wire	gpio6_4_zero,
	output wire	gpio6_4_one,
	output wire	gpio6_5_tie_hi_esd,
	input wire	[2:0]	gpio6_5_dm,
	input wire	gpio6_5_slow,
	input wire	gpio6_5_oe_n,
	output wire	gpio6_5_tie_lo_esd,
	input wire	gpio6_5_inp_dis,
	input wire	gpio6_5_enable_vddio,
	input wire	gpio6_5_vtrip_sel,
	input wire	[1:0]	gpio6_5_ib_mode_sel,
	input wire	gpio6_5_out,
	input wire	[1:0]	gpio6_5_slew_ctl,
	input wire	gpio6_5_analog_pol,
	input wire	gpio6_5_analog_sel,
	input wire	gpio6_5_hys_trim,
	input wire	gpio6_5_hld_ovr,
	output wire	gpio6_5_in_h,
	input wire	gpio6_5_enable_h,
	output wire	gpio6_5_in,
	input wire	gpio6_5_hld_h_n,
	input wire	gpio6_5_enable_vdda_h,
	input wire	gpio6_5_analog_en,
	input wire	gpio6_5_enable_inp_h,
	input wire	gpio6_5_enable_vswitch_h,
	inout wire	gpio6_5_pad_a_noesd_h,
	inout wire	gpio6_5_pad_a_esd_0_h,
	inout wire	gpio6_5_pad_a_esd_1_h,
	output wire	gpio6_5_zero,
	output wire	gpio6_5_one,
	output wire	gpio6_6_tie_hi_esd,
	input wire	[2:0]	gpio6_6_dm,
	input wire	gpio6_6_slow,
	input wire	gpio6_6_oe_n,
	output wire	gpio6_6_tie_lo_esd,
	input wire	gpio6_6_inp_dis,
	input wire	gpio6_6_enable_vddio,
	input wire	gpio6_6_vtrip_sel,
	input wire	[1:0]	gpio6_6_ib_mode_sel,
	input wire	gpio6_6_out,
	input wire	[1:0]	gpio6_6_slew_ctl,
	input wire	gpio6_6_analog_pol,
	input wire	gpio6_6_analog_sel,
	input wire	gpio6_6_hys_trim,
	input wire	gpio6_6_hld_ovr,
	output wire	gpio6_6_in_h,
	input wire	gpio6_6_enable_h,
	output wire	gpio6_6_in,
	input wire	gpio6_6_hld_h_n,
	input wire	gpio6_6_enable_vdda_h,
	input wire	gpio6_6_analog_en,
	input wire	gpio6_6_enable_inp_h,
	input wire	gpio6_6_enable_vswitch_h,
	inout wire	gpio6_6_pad_a_noesd_h,
	inout wire	gpio6_6_pad_a_esd_0_h,
	inout wire	gpio6_6_pad_a_esd_1_h,
	output wire	gpio6_6_zero,
	output wire	gpio6_6_one,
	output wire	gpio6_7_tie_hi_esd,
	input wire	[2:0]	gpio6_7_dm,
	input wire	gpio6_7_slow,
	input wire	gpio6_7_oe_n,
	output wire	gpio6_7_tie_lo_esd,
	input wire	gpio6_7_inp_dis,
	input wire	gpio6_7_enable_vddio,
	input wire	gpio6_7_vtrip_sel,
	input wire	[1:0]	gpio6_7_ib_mode_sel,
	input wire	gpio6_7_out,
	input wire	[1:0]	gpio6_7_slew_ctl,
	input wire	gpio6_7_analog_pol,
	input wire	gpio6_7_analog_sel,
	input wire	gpio6_7_hys_trim,
	input wire	gpio6_7_hld_ovr,
	output wire	gpio6_7_in_h,
	input wire	gpio6_7_enable_h,
	output wire	gpio6_7_in,
	input wire	gpio6_7_hld_h_n,
	input wire	gpio6_7_enable_vdda_h,
	input wire	gpio6_7_analog_en,
	input wire	gpio6_7_enable_inp_h,
	input wire	gpio6_7_enable_vswitch_h,
	inout wire	gpio6_7_pad_a_noesd_h,
	inout wire	gpio6_7_pad_a_esd_0_h,
	inout wire	gpio6_7_pad_a_esd_1_h,
	output wire	gpio6_7_zero,
	output wire	gpio6_7_one,
	output wire	gpio7_0_tie_lo_esd,
	output wire	gpio7_0_in,
	output wire	gpio7_0_tie_hi_esd,
	input wire	gpio7_0_enable_vddio,
	input wire	gpio7_0_slow,
	inout wire	gpio7_0_pad_a_esd_0_h,
	inout wire	gpio7_0_pad_a_esd_1_h,
	inout wire	gpio7_0_pad_a_noesd_h,
	input wire	gpio7_0_analog_en,
	input wire	gpio7_0_analog_pol,
	input wire	gpio7_0_inp_dis,
	input wire	gpio7_0_enable_inp_h,
	input wire	gpio7_0_enable_h,
	input wire	gpio7_0_hld_h_n,
	input wire	gpio7_0_analog_sel,
	input wire	[2:0]	gpio7_0_dm,
	input wire	gpio7_0_hld_ovr,
	input wire	gpio7_0_out,
	input wire	gpio7_0_enable_vswitch_h,
	input wire	gpio7_0_enable_vdda_h,
	input wire	gpio7_0_vtrip_sel,
	input wire	gpio7_0_ib_mode_sel,
	input wire	gpio7_0_oe_n,
	output wire	gpio7_0_in_h,
	output wire	gpio7_0_zero,
	output wire	gpio7_0_one,
	output wire	gpio7_1_tie_lo_esd,
	output wire	gpio7_1_in,
	output wire	gpio7_1_tie_hi_esd,
	input wire	gpio7_1_enable_vddio,
	input wire	gpio7_1_slow,
	inout wire	gpio7_1_pad_a_esd_0_h,
	inout wire	gpio7_1_pad_a_esd_1_h,
	inout wire	gpio7_1_pad_a_noesd_h,
	input wire	gpio7_1_analog_en,
	input wire	gpio7_1_analog_pol,
	input wire	gpio7_1_inp_dis,
	input wire	gpio7_1_enable_inp_h,
	input wire	gpio7_1_enable_h,
	input wire	gpio7_1_hld_h_n,
	input wire	gpio7_1_analog_sel,
	input wire	[2:0]	gpio7_1_dm,
	input wire	gpio7_1_hld_ovr,
	input wire	gpio7_1_out,
	input wire	gpio7_1_enable_vswitch_h,
	input wire	gpio7_1_enable_vdda_h,
	input wire	gpio7_1_vtrip_sel,
	input wire	gpio7_1_ib_mode_sel,
	input wire	gpio7_1_oe_n,
	output wire	gpio7_1_in_h,
	output wire	gpio7_1_zero,
	output wire	gpio7_1_one,
	output wire	gpio7_2_tie_lo_esd,
	output wire	gpio7_2_in,
	output wire	gpio7_2_tie_hi_esd,
	input wire	gpio7_2_enable_vddio,
	input wire	gpio7_2_slow,
	inout wire	gpio7_2_pad_a_esd_0_h,
	inout wire	gpio7_2_pad_a_esd_1_h,
	inout wire	gpio7_2_pad_a_noesd_h,
	input wire	gpio7_2_analog_en,
	input wire	gpio7_2_analog_pol,
	input wire	gpio7_2_inp_dis,
	input wire	gpio7_2_enable_inp_h,
	input wire	gpio7_2_enable_h,
	input wire	gpio7_2_hld_h_n,
	input wire	gpio7_2_analog_sel,
	input wire	[2:0]	gpio7_2_dm,
	input wire	gpio7_2_hld_ovr,
	input wire	gpio7_2_out,
	input wire	gpio7_2_enable_vswitch_h,
	input wire	gpio7_2_enable_vdda_h,
	input wire	gpio7_2_vtrip_sel,
	input wire	gpio7_2_ib_mode_sel,
	input wire	gpio7_2_oe_n,
	output wire	gpio7_2_in_h,
	output wire	gpio7_2_zero,
	output wire	gpio7_2_one,
	output wire	gpio7_3_tie_lo_esd,
	output wire	gpio7_3_in,
	output wire	gpio7_3_tie_hi_esd,
	input wire	gpio7_3_enable_vddio,
	input wire	gpio7_3_slow,
	inout wire	gpio7_3_pad_a_esd_0_h,
	inout wire	gpio7_3_pad_a_esd_1_h,
	inout wire	gpio7_3_pad_a_noesd_h,
	input wire	gpio7_3_analog_en,
	input wire	gpio7_3_analog_pol,
	input wire	gpio7_3_inp_dis,
	input wire	gpio7_3_enable_inp_h,
	input wire	gpio7_3_enable_h,
	input wire	gpio7_3_hld_h_n,
	input wire	gpio7_3_analog_sel,
	input wire	[2:0]	gpio7_3_dm,
	input wire	gpio7_3_hld_ovr,
	input wire	gpio7_3_out,
	input wire	gpio7_3_enable_vswitch_h,
	input wire	gpio7_3_enable_vdda_h,
	input wire	gpio7_3_vtrip_sel,
	input wire	gpio7_3_ib_mode_sel,
	input wire	gpio7_3_oe_n,
	output wire	gpio7_3_in_h,
	output wire	gpio7_3_zero,
	output wire	gpio7_3_one,
	output wire	gpio7_4_tie_lo_esd,
	output wire	gpio7_4_in,
	output wire	gpio7_4_tie_hi_esd,
	input wire	gpio7_4_enable_vddio,
	input wire	gpio7_4_slow,
	inout wire	gpio7_4_pad_a_esd_0_h,
	inout wire	gpio7_4_pad_a_esd_1_h,
	inout wire	gpio7_4_pad_a_noesd_h,
	input wire	gpio7_4_analog_en,
	input wire	gpio7_4_analog_pol,
	input wire	gpio7_4_inp_dis,
	input wire	gpio7_4_enable_inp_h,
	input wire	gpio7_4_enable_h,
	input wire	gpio7_4_hld_h_n,
	input wire	gpio7_4_analog_sel,
	input wire	[2:0]	gpio7_4_dm,
	input wire	gpio7_4_hld_ovr,
	input wire	gpio7_4_out,
	input wire	gpio7_4_enable_vswitch_h,
	input wire	gpio7_4_enable_vdda_h,
	input wire	gpio7_4_vtrip_sel,
	input wire	gpio7_4_ib_mode_sel,
	input wire	gpio7_4_oe_n,
	output wire	gpio7_4_in_h,
	output wire	gpio7_4_zero,
	output wire	gpio7_4_one,
	output wire	gpio7_5_tie_lo_esd,
	output wire	gpio7_5_in,
	output wire	gpio7_5_tie_hi_esd,
	input wire	gpio7_5_enable_vddio,
	input wire	gpio7_5_slow,
	inout wire	gpio7_5_pad_a_esd_0_h,
	inout wire	gpio7_5_pad_a_esd_1_h,
	inout wire	gpio7_5_pad_a_noesd_h,
	input wire	gpio7_5_analog_en,
	input wire	gpio7_5_analog_pol,
	input wire	gpio7_5_inp_dis,
	input wire	gpio7_5_enable_inp_h,
	input wire	gpio7_5_enable_h,
	input wire	gpio7_5_hld_h_n,
	input wire	gpio7_5_analog_sel,
	input wire	[2:0]	gpio7_5_dm,
	input wire	gpio7_5_hld_ovr,
	input wire	gpio7_5_out,
	input wire	gpio7_5_enable_vswitch_h,
	input wire	gpio7_5_enable_vdda_h,
	input wire	gpio7_5_vtrip_sel,
	input wire	gpio7_5_ib_mode_sel,
	input wire	gpio7_5_oe_n,
	output wire	gpio7_5_in_h,
	output wire	gpio7_5_zero,
	output wire	gpio7_5_one,
	output wire	gpio7_6_tie_lo_esd,
	output wire	gpio7_6_in,
	output wire	gpio7_6_tie_hi_esd,
	input wire	gpio7_6_enable_vddio,
	input wire	gpio7_6_slow,
	inout wire	gpio7_6_pad_a_esd_0_h,
	inout wire	gpio7_6_pad_a_esd_1_h,
	inout wire	gpio7_6_pad_a_noesd_h,
	input wire	gpio7_6_analog_en,
	input wire	gpio7_6_analog_pol,
	input wire	gpio7_6_inp_dis,
	input wire	gpio7_6_enable_inp_h,
	input wire	gpio7_6_enable_h,
	input wire	gpio7_6_hld_h_n,
	input wire	gpio7_6_analog_sel,
	input wire	[2:0]	gpio7_6_dm,
	input wire	gpio7_6_hld_ovr,
	input wire	gpio7_6_out,
	input wire	gpio7_6_enable_vswitch_h,
	input wire	gpio7_6_enable_vdda_h,
	input wire	gpio7_6_vtrip_sel,
	input wire	gpio7_6_ib_mode_sel,
	input wire	gpio7_6_oe_n,
	output wire	gpio7_6_in_h,
	output wire	gpio7_6_zero,
	output wire	gpio7_6_one,
	output wire	gpio7_7_tie_lo_esd,
	output wire	gpio7_7_in,
	output wire	gpio7_7_tie_hi_esd,
	input wire	gpio7_7_enable_vddio,
	input wire	gpio7_7_slow,
	inout wire	gpio7_7_pad_a_esd_0_h,
	inout wire	gpio7_7_pad_a_esd_1_h,
	inout wire	gpio7_7_pad_a_noesd_h,
	input wire	gpio7_7_analog_en,
	input wire	gpio7_7_analog_pol,
	input wire	gpio7_7_inp_dis,
	input wire	gpio7_7_enable_inp_h,
	input wire	gpio7_7_enable_h,
	input wire	gpio7_7_hld_h_n,
	input wire	gpio7_7_analog_sel,
	input wire	[2:0]	gpio7_7_dm,
	input wire	gpio7_7_hld_ovr,
	input wire	gpio7_7_out,
	input wire	gpio7_7_enable_vswitch_h,
	input wire	gpio7_7_enable_vdda_h,
	input wire	gpio7_7_vtrip_sel,
	input wire	gpio7_7_ib_mode_sel,
	input wire	gpio7_7_oe_n,
	output wire	gpio7_7_in_h,
	output wire	gpio7_7_zero,
	output wire	gpio7_7_one,
	input wire	muxsplit_sw_hld_vdda_h_n,
	input wire	muxsplit_sw_enable_vdda_h,
	input wire	muxsplit_sw_switch_aa_sl,
	input wire	muxsplit_sw_switch_aa_s0,
	input wire	muxsplit_sw_switch_bb_s0,
	input wire	muxsplit_sw_switch_bb_sl,
	input wire	muxsplit_sw_switch_bb_sr,
	input wire	muxsplit_sw_switch_aa_sr
);

	/* Declaration of wires internal to the padframe and not connected
	 * to a padframe pin.
	 */

	wire amuxbus_a_e;
	wire amuxbus_b_e;
	wire amuxbus_a_w;
	wire amuxbus_b_w;
	wire amuxbus_a_s;
	wire amuxbus_b_s;

	wire vddio_q;
	wire vssio_q;
	
    sky130_fd_io__top_gpio_ovtv2 gpio1_0_pad (
	.OUT(gpio1_0_out),
	.OE_N(gpio1_0_oe_n),
	.HLD_H_N(gpio1_0_hld_h_n),
	.ENABLE_H(gpio1_0_enable_h),
	.ENABLE_INP_H(gpio1_0_enable_inp_h),
	.ENABLE_VDDA_H(gpio1_0_enable_vdda_h),
	.ENABLE_VDDIO(gpio1_0_enable_vddio),
	.ENABLE_VSWITCH_H(gpio1_0_enable_vswitch_h),
	.INP_DIS(gpio1_0_inp_dis),
	.VTRIP_SEL(gpio1_0_vtrip_sel),
	.HYS_TRIM(gpio1_0_hys_trim),
	.SLOW(gpio1_0_slow),
	.SLEW_CTL(gpio1_0_slew_ctl),
	.HLD_OVR(gpio1_0_hld_ovr),
	.ANALOG_EN(gpio1_0_analog_en),
	.ANALOG_SEL(gpio1_0_analog_sel),
	.ANALOG_POL(gpio1_0_analog_pol),
	.DM(gpio1_0_dm),
	.IB_MODE_SEL(gpio1_0_ib_mode_sel),
	.VINREF(vref_e_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda1),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio1_0),
	.PAD_A_NOESD_H(gpio1_0_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio1_0_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio1_0_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.IN(gpio1_0_in),
	.IN_H(gpio1_0_in_h),
	.TIE_HI_ESD(gpio1_0_tie_hi_esd),
	.TIE_LO_ESD(gpio1_0_tie_lo_esd)
    );

    constant_block gpio1_0_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio1_0_one),
	.zero(gpio1_0_zero)
    );

    sky130_ef_io__gpiov2_pad gpio3_3_pad (
	.IN_H(gpio3_3_in_h),
	.IN(gpio3_3_in),
	.OUT(gpio3_3_out),
	.OE_N(gpio3_3_oe_n),
	.HLD_H_N(gpio3_3_hld_h_n),
	.ENABLE_H(gpio3_3_enable_h),
	.ENABLE_INP_H(gpio3_3_enable_inp_h),
	.ENABLE_VDDA_H(gpio3_3_enable_vdda_h),
	.ENABLE_VDDIO(gpio3_3_enable_vddio),
	.ENABLE_VSWITCH_H(gpio3_3_enable_vswitch_h),
	.INP_DIS(gpio3_3_inp_dis),
	.VTRIP_SEL(gpio3_3_vtrip_sel),
	.SLOW(gpio3_3_slow),
	.HLD_OVR(gpio3_3_hld_ovr),
	.ANALOG_EN(gpio3_3_analog_en),
	.ANALOG_SEL(gpio3_3_analog_sel),
	.ANALOG_POL(gpio3_3_analog_pol),
	.DM(gpio3_3_dm),
	.IB_MODE_SEL(gpio3_3_ib_mode_sel),
	.PAD(gpio3_3),
	.PAD_A_NOESD_H(gpio3_3_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio3_3_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio3_3_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio3_3_tie_hi_esd),
	.TIE_LO_ESD(gpio3_3_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio3_3_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio3_3_one),
	.zero(gpio3_3_zero)
    );

    sky130_ef_io__vssio_hvc_clamped_pad vssio_2_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VSSIO_PAD(vssio_2),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio5_6_pad (
	.IN_H(gpio5_6_in_h),
	.IN(gpio5_6_in),
	.OUT(gpio5_6_out),
	.OE_N(gpio5_6_oe_n),
	.HLD_H_N(gpio5_6_hld_h_n),
	.ENABLE_H(gpio5_6_enable_h),
	.ENABLE_INP_H(gpio5_6_enable_inp_h),
	.ENABLE_VDDA_H(gpio5_6_enable_vdda_h),
	.ENABLE_VDDIO(gpio5_6_enable_vddio),
	.ENABLE_VSWITCH_H(gpio5_6_enable_vswitch_h),
	.INP_DIS(gpio5_6_inp_dis),
	.VTRIP_SEL(gpio5_6_vtrip_sel),
	.SLOW(gpio5_6_slow),
	.HLD_OVR(gpio5_6_hld_ovr),
	.ANALOG_EN(gpio5_6_analog_en),
	.ANALOG_SEL(gpio5_6_analog_sel),
	.ANALOG_POL(gpio5_6_analog_pol),
	.DM(gpio5_6_dm),
	.IB_MODE_SEL(gpio5_6_ib_mode_sel),
	.PAD(gpio5_6),
	.PAD_A_NOESD_H(gpio5_6_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio5_6_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio5_6_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio5_6_tie_hi_esd),
	.TIE_LO_ESD(gpio5_6_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio5_6_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio5_6_one),
	.zero(gpio5_6_zero)
    );

    sky130_ef_io__vddio_hvc_clamped_pad vddio_3_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VDDIO_PAD(vddio_3),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio0_0_pad (
	.IN_H(gpio0_0_in_h),
	.IN(gpio0_0_in),
	.OUT(gpio0_0_out),
	.OE_N(gpio0_0_oe_n),
	.HLD_H_N(gpio0_0_hld_h_n),
	.ENABLE_H(gpio0_0_enable_h),
	.ENABLE_INP_H(gpio0_0_enable_inp_h),
	.ENABLE_VDDA_H(gpio0_0_enable_vdda_h),
	.ENABLE_VDDIO(gpio0_0_enable_vddio),
	.ENABLE_VSWITCH_H(gpio0_0_enable_vswitch_h),
	.INP_DIS(gpio0_0_inp_dis),
	.VTRIP_SEL(gpio0_0_vtrip_sel),
	.SLOW(gpio0_0_slow),
	.HLD_OVR(gpio0_0_hld_ovr),
	.ANALOG_EN(gpio0_0_analog_en),
	.ANALOG_SEL(gpio0_0_analog_sel),
	.ANALOG_POL(gpio0_0_analog_pol),
	.DM(gpio0_0_dm),
	.IB_MODE_SEL(gpio0_0_ib_mode_sel),
	.PAD(gpio0_0),
	.PAD_A_NOESD_H(gpio0_0_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio0_0_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio0_0_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio0_0_tie_hi_esd),
	.TIE_LO_ESD(gpio0_0_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio0_0_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio0_0_one),
	.zero(gpio0_0_zero)
    );

    sky130_ef_io__gpiov2_pad gpio2_3_pad (
	.IN_H(gpio2_3_in_h),
	.IN(gpio2_3_in),
	.OUT(gpio2_3_out),
	.OE_N(gpio2_3_oe_n),
	.HLD_H_N(gpio2_3_hld_h_n),
	.ENABLE_H(gpio2_3_enable_h),
	.ENABLE_INP_H(gpio2_3_enable_inp_h),
	.ENABLE_VDDA_H(gpio2_3_enable_vdda_h),
	.ENABLE_VDDIO(gpio2_3_enable_vddio),
	.ENABLE_VSWITCH_H(gpio2_3_enable_vswitch_h),
	.INP_DIS(gpio2_3_inp_dis),
	.VTRIP_SEL(gpio2_3_vtrip_sel),
	.SLOW(gpio2_3_slow),
	.HLD_OVR(gpio2_3_hld_ovr),
	.ANALOG_EN(gpio2_3_analog_en),
	.ANALOG_SEL(gpio2_3_analog_sel),
	.ANALOG_POL(gpio2_3_analog_pol),
	.DM(gpio2_3_dm),
	.IB_MODE_SEL(gpio2_3_ib_mode_sel),
	.PAD(gpio2_3),
	.PAD_A_NOESD_H(gpio2_3_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio2_3_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio2_3_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio2_3_tie_hi_esd),
	.TIE_LO_ESD(gpio2_3_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio2_3_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio2_3_one),
	.zero(gpio2_3_zero)
    );

    sky130_ef_io__gpiov2_pad gpio4_6_pad (
	.IN_H(gpio4_6_in_h),
	.IN(gpio4_6_in),
	.OUT(gpio4_6_out),
	.OE_N(gpio4_6_oe_n),
	.HLD_H_N(gpio4_6_hld_h_n),
	.ENABLE_H(gpio4_6_enable_h),
	.ENABLE_INP_H(gpio4_6_enable_inp_h),
	.ENABLE_VDDA_H(gpio4_6_enable_vdda_h),
	.ENABLE_VDDIO(gpio4_6_enable_vddio),
	.ENABLE_VSWITCH_H(gpio4_6_enable_vswitch_h),
	.INP_DIS(gpio4_6_inp_dis),
	.VTRIP_SEL(gpio4_6_vtrip_sel),
	.SLOW(gpio4_6_slow),
	.HLD_OVR(gpio4_6_hld_ovr),
	.ANALOG_EN(gpio4_6_analog_en),
	.ANALOG_SEL(gpio4_6_analog_sel),
	.ANALOG_POL(gpio4_6_analog_pol),
	.DM(gpio4_6_dm),
	.IB_MODE_SEL(gpio4_6_ib_mode_sel),
	.PAD(gpio4_6),
	.PAD_A_NOESD_H(gpio4_6_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio4_6_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio4_6_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio4_6_tie_hi_esd),
	.TIE_LO_ESD(gpio4_6_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio4_6_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio4_6_one),
	.zero(gpio4_6_zero)
    );

    sky130_fd_io__top_gpiovrefv2 vref_w (
	.amuxbus_a(amuxbus_a_w),
	.amuxbus_b(amuxbus_b_w),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda2),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa2),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio),
	.enable_h(vref_w_enable_h),
	.hld_h_n(vref_w_hld_h_n),
	.ref_sel(vref_w_ref_sel),
	.vrefgen_en(vref_w_vrefgen_en),
	.vinref(vref_w_vinref)
    );

    sky130_ef_io__vssa_hvc_clamped_pad vssa2_1_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VSSA_PAD(vssa2_1),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_fd_io__top_gpio_ovtv2 gpio1_3_pad (
	.OUT(gpio1_3_out),
	.OE_N(gpio1_3_oe_n),
	.HLD_H_N(gpio1_3_hld_h_n),
	.ENABLE_H(gpio1_3_enable_h),
	.ENABLE_INP_H(gpio1_3_enable_inp_h),
	.ENABLE_VDDA_H(gpio1_3_enable_vdda_h),
	.ENABLE_VDDIO(gpio1_3_enable_vddio),
	.ENABLE_VSWITCH_H(gpio1_3_enable_vswitch_h),
	.INP_DIS(gpio1_3_inp_dis),
	.VTRIP_SEL(gpio1_3_vtrip_sel),
	.HYS_TRIM(gpio1_3_hys_trim),
	.SLOW(gpio1_3_slow),
	.SLEW_CTL(gpio1_3_slew_ctl),
	.HLD_OVR(gpio1_3_hld_ovr),
	.ANALOG_EN(gpio1_3_analog_en),
	.ANALOG_SEL(gpio1_3_analog_sel),
	.ANALOG_POL(gpio1_3_analog_pol),
	.DM(gpio1_3_dm),
	.IB_MODE_SEL(gpio1_3_ib_mode_sel),
	.VINREF(vref_e_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda1),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio1_3),
	.PAD_A_NOESD_H(gpio1_3_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio1_3_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio1_3_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.IN(gpio1_3_in),
	.IN_H(gpio1_3_in_h),
	.TIE_HI_ESD(gpio1_3_tie_hi_esd),
	.TIE_LO_ESD(gpio1_3_tie_lo_esd)
    );

    constant_block gpio1_3_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio1_3_one),
	.zero(gpio1_3_zero)
    );

    sky130_ef_io__vssio_hvc_clamped_pad vssio_5_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VSSIO_PAD(vssio_5),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio3_6_pad (
	.IN_H(gpio3_6_in_h),
	.IN(gpio3_6_in),
	.OUT(gpio3_6_out),
	.OE_N(gpio3_6_oe_n),
	.HLD_H_N(gpio3_6_hld_h_n),
	.ENABLE_H(gpio3_6_enable_h),
	.ENABLE_INP_H(gpio3_6_enable_inp_h),
	.ENABLE_VDDA_H(gpio3_6_enable_vdda_h),
	.ENABLE_VDDIO(gpio3_6_enable_vddio),
	.ENABLE_VSWITCH_H(gpio3_6_enable_vswitch_h),
	.INP_DIS(gpio3_6_inp_dis),
	.VTRIP_SEL(gpio3_6_vtrip_sel),
	.SLOW(gpio3_6_slow),
	.HLD_OVR(gpio3_6_hld_ovr),
	.ANALOG_EN(gpio3_6_analog_en),
	.ANALOG_SEL(gpio3_6_analog_sel),
	.ANALOG_POL(gpio3_6_analog_pol),
	.DM(gpio3_6_dm),
	.IB_MODE_SEL(gpio3_6_ib_mode_sel),
	.PAD(gpio3_6),
	.PAD_A_NOESD_H(gpio3_6_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio3_6_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio3_6_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio3_6_tie_hi_esd),
	.TIE_LO_ESD(gpio3_6_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio3_6_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio3_6_one),
	.zero(gpio3_6_zero)
    );

    sky130_fd_io__top_amuxsplitv2 muxsplit_se (
	.amuxbus_a_l(amuxbus_a_e),
	.amuxbus_a_r(amuxbus_a_s),
	.amuxbus_b_l(amuxbus_b_e),
	.amuxbus_b_r(amuxbus_b_s),
	.enable_vdda_h(muxsplit_se_enable_vdda_h),
	.hld_vdda_h_n(muxsplit_se_hld_vdda_h_n),
	.switch_aa_s0(muxsplit_se_switch_aa_s0),
	.switch_aa_sl(muxsplit_se_switch_aa_sl),
	.switch_aa_sr(muxsplit_se_switch_aa_sr),
	.switch_bb_s0(muxsplit_se_switch_bb_s0),
	.switch_bb_sl(muxsplit_se_switch_bb_sl),
	.switch_bb_sr(muxsplit_se_switch_bb_sr),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda3),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa3),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio)
    );

    sky130_ef_io__vssa_hvc_clamped_pad vssa1_1_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VSSA_PAD(vssa1_1),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__vddio_hvc_clamped_pad vddio_6_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VDDIO_PAD(vddio_6),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio0_3_pad (
	.IN_H(gpio0_3_in_h),
	.IN(gpio0_3_in),
	.OUT(gpio0_3_out),
	.OE_N(gpio0_3_oe_n),
	.HLD_H_N(gpio0_3_hld_h_n),
	.ENABLE_H(gpio0_3_enable_h),
	.ENABLE_INP_H(gpio0_3_enable_inp_h),
	.ENABLE_VDDA_H(gpio0_3_enable_vdda_h),
	.ENABLE_VDDIO(gpio0_3_enable_vddio),
	.ENABLE_VSWITCH_H(gpio0_3_enable_vswitch_h),
	.INP_DIS(gpio0_3_inp_dis),
	.VTRIP_SEL(gpio0_3_vtrip_sel),
	.SLOW(gpio0_3_slow),
	.HLD_OVR(gpio0_3_hld_ovr),
	.ANALOG_EN(gpio0_3_analog_en),
	.ANALOG_SEL(gpio0_3_analog_sel),
	.ANALOG_POL(gpio0_3_analog_pol),
	.DM(gpio0_3_dm),
	.IB_MODE_SEL(gpio0_3_ib_mode_sel),
	.PAD(gpio0_3),
	.PAD_A_NOESD_H(gpio0_3_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio0_3_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio0_3_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio0_3_tie_hi_esd),
	.TIE_LO_ESD(gpio0_3_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio0_3_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio0_3_one),
	.zero(gpio0_3_zero)
    );

    sky130_ef_io__gpiov2_pad gpio2_6_pad (
	.IN_H(gpio2_6_in_h),
	.IN(gpio2_6_in),
	.OUT(gpio2_6_out),
	.OE_N(gpio2_6_oe_n),
	.HLD_H_N(gpio2_6_hld_h_n),
	.ENABLE_H(gpio2_6_enable_h),
	.ENABLE_INP_H(gpio2_6_enable_inp_h),
	.ENABLE_VDDA_H(gpio2_6_enable_vdda_h),
	.ENABLE_VDDIO(gpio2_6_enable_vddio),
	.ENABLE_VSWITCH_H(gpio2_6_enable_vswitch_h),
	.INP_DIS(gpio2_6_inp_dis),
	.VTRIP_SEL(gpio2_6_vtrip_sel),
	.SLOW(gpio2_6_slow),
	.HLD_OVR(gpio2_6_hld_ovr),
	.ANALOG_EN(gpio2_6_analog_en),
	.ANALOG_SEL(gpio2_6_analog_sel),
	.ANALOG_POL(gpio2_6_analog_pol),
	.DM(gpio2_6_dm),
	.IB_MODE_SEL(gpio2_6_ib_mode_sel),
	.PAD(gpio2_6),
	.PAD_A_NOESD_H(gpio2_6_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio2_6_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio2_6_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio2_6_tie_hi_esd),
	.TIE_LO_ESD(gpio2_6_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio2_6_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio2_6_one),
	.zero(gpio2_6_zero)
    );

    sky130_fd_io__top_analog_pad xo0_pad (
	.pad_core(xo0_core),
	.pad(xo0),
	.amuxbus_a(amuxbus_a_s),
	.amuxbus_b(amuxbus_b_s),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda3),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa3),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio8_2_pad (
	.IN_H(gpio8_2_in_h),
	.IN(gpio8_2_in),
	.OUT(gpio8_2_out),
	.OE_N(gpio8_2_oe_n),
	.HLD_H_N(gpio8_2_hld_h_n),
	.ENABLE_H(gpio8_2_enable_h),
	.ENABLE_INP_H(gpio8_2_enable_inp_h),
	.ENABLE_VDDA_H(gpio8_2_enable_vdda_h),
	.ENABLE_VDDIO(gpio8_2_enable_vddio),
	.ENABLE_VSWITCH_H(gpio8_2_enable_vswitch_h),
	.INP_DIS(gpio8_2_inp_dis),
	.VTRIP_SEL(gpio8_2_vtrip_sel),
	.SLOW(gpio8_2_slow),
	.HLD_OVR(gpio8_2_hld_ovr),
	.ANALOG_EN(gpio8_2_analog_en),
	.ANALOG_SEL(gpio8_2_analog_sel),
	.ANALOG_POL(gpio8_2_analog_pol),
	.DM(gpio8_2_dm),
	.IB_MODE_SEL(gpio8_2_ib_mode_sel),
	.PAD(gpio8_2),
	.PAD_A_NOESD_H(gpio8_2_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio8_2_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio8_2_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio8_2_tie_hi_esd),
	.TIE_LO_ESD(gpio8_2_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio8_2_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio8_2_one),
	.zero(gpio8_2_zero)
    );

    sky130_fd_io__top_gpio_ovtv2 gpio1_6_pad (
	.OUT(gpio1_6_out),
	.OE_N(gpio1_6_oe_n),
	.HLD_H_N(gpio1_6_hld_h_n),
	.ENABLE_H(gpio1_6_enable_h),
	.ENABLE_INP_H(gpio1_6_enable_inp_h),
	.ENABLE_VDDA_H(gpio1_6_enable_vdda_h),
	.ENABLE_VDDIO(gpio1_6_enable_vddio),
	.ENABLE_VSWITCH_H(gpio1_6_enable_vswitch_h),
	.INP_DIS(gpio1_6_inp_dis),
	.VTRIP_SEL(gpio1_6_vtrip_sel),
	.HYS_TRIM(gpio1_6_hys_trim),
	.SLOW(gpio1_6_slow),
	.SLEW_CTL(gpio1_6_slew_ctl),
	.HLD_OVR(gpio1_6_hld_ovr),
	.ANALOG_EN(gpio1_6_analog_en),
	.ANALOG_SEL(gpio1_6_analog_sel),
	.ANALOG_POL(gpio1_6_analog_pol),
	.DM(gpio1_6_dm),
	.IB_MODE_SEL(gpio1_6_ib_mode_sel),
	.VINREF(vref_e_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda1),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio1_6),
	.PAD_A_NOESD_H(gpio1_6_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio1_6_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio1_6_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.IN(gpio1_6_in),
	.IN_H(gpio1_6_in_h),
	.TIE_HI_ESD(gpio1_6_tie_hi_esd),
	.TIE_LO_ESD(gpio1_6_tie_lo_esd)
    );

    constant_block gpio1_6_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio1_6_one),
	.zero(gpio1_6_zero)
    );

    sky130_ef_io__vssio_hvc_clamped_pad vssio_8_pad (
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VSSIO_PAD(vssio_8),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__vccd_lvc_clamped3_pad vccd2_2_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD_PAD(vccd2_2),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio),
	.VCCD1(vccd2[5]),
	.VSSD1(vssd2[5])
    );

    sky130_ef_io__gpiov2_pad gpio7_2_pad (
	.IN_H(gpio7_2_in_h),
	.IN(gpio7_2_in),
	.OUT(gpio7_2_out),
	.OE_N(gpio7_2_oe_n),
	.HLD_H_N(gpio7_2_hld_h_n),
	.ENABLE_H(gpio7_2_enable_h),
	.ENABLE_INP_H(gpio7_2_enable_inp_h),
	.ENABLE_VDDA_H(gpio7_2_enable_vdda_h),
	.ENABLE_VDDIO(gpio7_2_enable_vddio),
	.ENABLE_VSWITCH_H(gpio7_2_enable_vswitch_h),
	.INP_DIS(gpio7_2_inp_dis),
	.VTRIP_SEL(gpio7_2_vtrip_sel),
	.SLOW(gpio7_2_slow),
	.HLD_OVR(gpio7_2_hld_ovr),
	.ANALOG_EN(gpio7_2_analog_en),
	.ANALOG_SEL(gpio7_2_analog_sel),
	.ANALOG_POL(gpio7_2_analog_pol),
	.DM(gpio7_2_dm),
	.IB_MODE_SEL(gpio7_2_ib_mode_sel),
	.PAD(gpio7_2),
	.PAD_A_NOESD_H(gpio7_2_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio7_2_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio7_2_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio7_2_tie_hi_esd),
	.TIE_LO_ESD(gpio7_2_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio7_2_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio7_2_one),
	.zero(gpio7_2_zero)
    );

    sky130_ef_io__vddio_hvc_clamped_pad vddio_9_pad (
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VCCD(vccd0),
	.VDDIO_PAD(vddio_9),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio0_6_pad (
	.IN_H(gpio0_6_in_h),
	.IN(gpio0_6_in),
	.OUT(gpio0_6_out),
	.OE_N(gpio0_6_oe_n),
	.HLD_H_N(gpio0_6_hld_h_n),
	.ENABLE_H(gpio0_6_enable_h),
	.ENABLE_INP_H(gpio0_6_enable_inp_h),
	.ENABLE_VDDA_H(gpio0_6_enable_vdda_h),
	.ENABLE_VDDIO(gpio0_6_enable_vddio),
	.ENABLE_VSWITCH_H(gpio0_6_enable_vswitch_h),
	.INP_DIS(gpio0_6_inp_dis),
	.VTRIP_SEL(gpio0_6_vtrip_sel),
	.SLOW(gpio0_6_slow),
	.HLD_OVR(gpio0_6_hld_ovr),
	.ANALOG_EN(gpio0_6_analog_en),
	.ANALOG_SEL(gpio0_6_analog_sel),
	.ANALOG_POL(gpio0_6_analog_pol),
	.DM(gpio0_6_dm),
	.IB_MODE_SEL(gpio0_6_ib_mode_sel),
	.PAD(gpio0_6),
	.PAD_A_NOESD_H(gpio0_6_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio0_6_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio0_6_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio0_6_tie_hi_esd),
	.TIE_LO_ESD(gpio0_6_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio0_6_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio0_6_one),
	.zero(gpio0_6_zero)
    );

    sky130_ef_io__vccd_lvc_clamped3_pad vccd1_2_pad (
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD_PAD(vccd1_2),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio),
	.VCCD1(vccd1[5]),
	.VSSD1(vssd1[5])
    );

    sky130_fd_io__top_gpio_ovtv2 gpio6_2_pad (
	.OUT(gpio6_2_out),
	.OE_N(gpio6_2_oe_n),
	.HLD_H_N(gpio6_2_hld_h_n),
	.ENABLE_H(gpio6_2_enable_h),
	.ENABLE_INP_H(gpio6_2_enable_inp_h),
	.ENABLE_VDDA_H(gpio6_2_enable_vdda_h),
	.ENABLE_VDDIO(gpio6_2_enable_vddio),
	.ENABLE_VSWITCH_H(gpio6_2_enable_vswitch_h),
	.INP_DIS(gpio6_2_inp_dis),
	.VTRIP_SEL(gpio6_2_vtrip_sel),
	.HYS_TRIM(gpio6_2_hys_trim),
	.SLOW(gpio6_2_slow),
	.SLEW_CTL(gpio6_2_slew_ctl),
	.HLD_OVR(gpio6_2_hld_ovr),
	.ANALOG_EN(gpio6_2_analog_en),
	.ANALOG_SEL(gpio6_2_analog_sel),
	.ANALOG_POL(gpio6_2_analog_pol),
	.DM(gpio6_2_dm),
	.IB_MODE_SEL(gpio6_2_ib_mode_sel),
	.VINREF(vref_e_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda2),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio6_2),
	.PAD_A_NOESD_H(gpio6_2_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio6_2_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio6_2_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.IN(gpio6_2_in),
	.IN_H(gpio6_2_in_h),
	.TIE_HI_ESD(gpio6_2_tie_hi_esd),
	.TIE_LO_ESD(gpio6_2_tie_lo_esd)
    );

    constant_block gpio6_2_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio6_2_one),
	.zero(gpio6_2_zero)
    );

    sky130_ef_io__gpiov2_pad gpio8_5_pad (
	.IN_H(gpio8_5_in_h),
	.IN(gpio8_5_in),
	.OUT(gpio8_5_out),
	.OE_N(gpio8_5_oe_n),
	.HLD_H_N(gpio8_5_hld_h_n),
	.ENABLE_H(gpio8_5_enable_h),
	.ENABLE_INP_H(gpio8_5_enable_inp_h),
	.ENABLE_VDDA_H(gpio8_5_enable_vdda_h),
	.ENABLE_VDDIO(gpio8_5_enable_vddio),
	.ENABLE_VSWITCH_H(gpio8_5_enable_vswitch_h),
	.INP_DIS(gpio8_5_inp_dis),
	.VTRIP_SEL(gpio8_5_vtrip_sel),
	.SLOW(gpio8_5_slow),
	.HLD_OVR(gpio8_5_hld_ovr),
	.ANALOG_EN(gpio8_5_analog_en),
	.ANALOG_SEL(gpio8_5_analog_sel),
	.ANALOG_POL(gpio8_5_analog_pol),
	.DM(gpio8_5_dm),
	.IB_MODE_SEL(gpio8_5_ib_mode_sel),
	.PAD(gpio8_5),
	.PAD_A_NOESD_H(gpio8_5_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio8_5_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio8_5_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio8_5_tie_hi_esd),
	.TIE_LO_ESD(gpio8_5_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio8_5_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio8_5_one),
	.zero(gpio8_5_zero)
    );

    sky130_fd_io__top_amuxsplitv2 muxsplit_ne (
	.amuxbus_a_l(amuxbus_a_n),
	.amuxbus_a_r(amuxbus_a_e),
	.amuxbus_b_l(amuxbus_b_n),
	.amuxbus_b_r(amuxbus_b_e),
	.enable_vdda_h(muxsplit_ne_enable_vdda_h),
	.hld_vdda_h_n(muxsplit_ne_hld_vdda_h_n),
	.switch_aa_s0(muxsplit_ne_switch_aa_s0),
	.switch_aa_sl(muxsplit_ne_switch_aa_sl),
	.switch_aa_sr(muxsplit_ne_switch_aa_sr),
	.switch_bb_s0(muxsplit_ne_switch_bb_s0),
	.switch_bb_sl(muxsplit_ne_switch_bb_sl),
	.switch_bb_sr(muxsplit_ne_switch_bb_sr),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda0),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa0),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio5_2_pad (
	.IN_H(gpio5_2_in_h),
	.IN(gpio5_2_in),
	.OUT(gpio5_2_out),
	.OE_N(gpio5_2_oe_n),
	.HLD_H_N(gpio5_2_hld_h_n),
	.ENABLE_H(gpio5_2_enable_h),
	.ENABLE_INP_H(gpio5_2_enable_inp_h),
	.ENABLE_VDDA_H(gpio5_2_enable_vdda_h),
	.ENABLE_VDDIO(gpio5_2_enable_vddio),
	.ENABLE_VSWITCH_H(gpio5_2_enable_vswitch_h),
	.INP_DIS(gpio5_2_inp_dis),
	.VTRIP_SEL(gpio5_2_vtrip_sel),
	.SLOW(gpio5_2_slow),
	.HLD_OVR(gpio5_2_hld_ovr),
	.ANALOG_EN(gpio5_2_analog_en),
	.ANALOG_SEL(gpio5_2_analog_sel),
	.ANALOG_POL(gpio5_2_analog_pol),
	.DM(gpio5_2_dm),
	.IB_MODE_SEL(gpio5_2_ib_mode_sel),
	.PAD(gpio5_2),
	.PAD_A_NOESD_H(gpio5_2_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio5_2_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio5_2_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio5_2_tie_hi_esd),
	.TIE_LO_ESD(gpio5_2_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio5_2_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio5_2_one),
	.zero(gpio5_2_zero)
    );

    sky130_ef_io__gpiov2_pad gpio7_5_pad (
	.IN_H(gpio7_5_in_h),
	.IN(gpio7_5_in),
	.OUT(gpio7_5_out),
	.OE_N(gpio7_5_oe_n),
	.HLD_H_N(gpio7_5_hld_h_n),
	.ENABLE_H(gpio7_5_enable_h),
	.ENABLE_INP_H(gpio7_5_enable_inp_h),
	.ENABLE_VDDA_H(gpio7_5_enable_vdda_h),
	.ENABLE_VDDIO(gpio7_5_enable_vddio),
	.ENABLE_VSWITCH_H(gpio7_5_enable_vswitch_h),
	.INP_DIS(gpio7_5_inp_dis),
	.VTRIP_SEL(gpio7_5_vtrip_sel),
	.SLOW(gpio7_5_slow),
	.HLD_OVR(gpio7_5_hld_ovr),
	.ANALOG_EN(gpio7_5_analog_en),
	.ANALOG_SEL(gpio7_5_analog_sel),
	.ANALOG_POL(gpio7_5_analog_pol),
	.DM(gpio7_5_dm),
	.IB_MODE_SEL(gpio7_5_ib_mode_sel),
	.PAD(gpio7_5),
	.PAD_A_NOESD_H(gpio7_5_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio7_5_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio7_5_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio7_5_tie_hi_esd),
	.TIE_LO_ESD(gpio7_5_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio7_5_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio7_5_one),
	.zero(gpio7_5_zero)
    );

    sky130_fd_io__top_analog_pad analog_0_pad (
	.pad_core(analog_0_core),
	.pad(analog_0),
	.amuxbus_a(amuxbus_a_n),
	.amuxbus_b(amuxbus_b_n),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda0),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa0),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio4_2_pad (
	.IN_H(gpio4_2_in_h),
	.IN(gpio4_2_in),
	.OUT(gpio4_2_out),
	.OE_N(gpio4_2_oe_n),
	.HLD_H_N(gpio4_2_hld_h_n),
	.ENABLE_H(gpio4_2_enable_h),
	.ENABLE_INP_H(gpio4_2_enable_inp_h),
	.ENABLE_VDDA_H(gpio4_2_enable_vdda_h),
	.ENABLE_VDDIO(gpio4_2_enable_vddio),
	.ENABLE_VSWITCH_H(gpio4_2_enable_vswitch_h),
	.INP_DIS(gpio4_2_inp_dis),
	.VTRIP_SEL(gpio4_2_vtrip_sel),
	.SLOW(gpio4_2_slow),
	.HLD_OVR(gpio4_2_hld_ovr),
	.ANALOG_EN(gpio4_2_analog_en),
	.ANALOG_SEL(gpio4_2_analog_sel),
	.ANALOG_POL(gpio4_2_analog_pol),
	.DM(gpio4_2_dm),
	.IB_MODE_SEL(gpio4_2_ib_mode_sel),
	.PAD(gpio4_2),
	.PAD_A_NOESD_H(gpio4_2_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio4_2_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio4_2_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio4_2_tie_hi_esd),
	.TIE_LO_ESD(gpio4_2_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio4_2_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio4_2_one),
	.zero(gpio4_2_zero)
    );

    sky130_ef_io__vssd_lvc_clamped3_pad vssd2_2_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VSSD_PAD(vssd2_2),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio),
	.VCCD1(vccd2[4]),
	.VSSD1(vssd2[4])
    );

    sky130_fd_io__top_gpio_ovtv2 gpio6_5_pad (
	.OUT(gpio6_5_out),
	.OE_N(gpio6_5_oe_n),
	.HLD_H_N(gpio6_5_hld_h_n),
	.ENABLE_H(gpio6_5_enable_h),
	.ENABLE_INP_H(gpio6_5_enable_inp_h),
	.ENABLE_VDDA_H(gpio6_5_enable_vdda_h),
	.ENABLE_VDDIO(gpio6_5_enable_vddio),
	.ENABLE_VSWITCH_H(gpio6_5_enable_vswitch_h),
	.INP_DIS(gpio6_5_inp_dis),
	.VTRIP_SEL(gpio6_5_vtrip_sel),
	.HYS_TRIM(gpio6_5_hys_trim),
	.SLOW(gpio6_5_slow),
	.SLEW_CTL(gpio6_5_slew_ctl),
	.HLD_OVR(gpio6_5_hld_ovr),
	.ANALOG_EN(gpio6_5_analog_en),
	.ANALOG_SEL(gpio6_5_analog_sel),
	.ANALOG_POL(gpio6_5_analog_pol),
	.DM(gpio6_5_dm),
	.IB_MODE_SEL(gpio6_5_ib_mode_sel),
	.VINREF(vref_w_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda2),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio6_5),
	.PAD_A_NOESD_H(gpio6_5_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio6_5_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio6_5_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.IN(gpio6_5_in),
	.IN_H(gpio6_5_in_h),
	.TIE_HI_ESD(gpio6_5_tie_hi_esd),
	.TIE_LO_ESD(gpio6_5_tie_lo_esd)
    );

    constant_block gpio6_5_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio6_5_one),
	.zero(gpio6_5_zero)
    );

    sky130_fd_io__top_sio_macro sio_macro_pads (
	.OUT(sio_out),
	.OE_N(sio_oe_n),
	.HLD_H_N(sio_hld_h_n),
	.ENABLE_H(sio_enable_h),
	.ENABLE_VDDA_H(sio_enable_vdda_h),
	.INP_DIS(sio_inp_dis),
	.VTRIP_SEL(sio_vtrip_sel),
	.SLOW(sio_slow),
	.HLD_OVR(sio_hld_ovr),
	.IBUF_SEL(sio_ibuf_sel),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda3),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD({sio0, sio1}),
	.PAD_A_NOESD_H(sio_pad_a_noesd_h),
	.PAD_A_ESD_0_H(sio_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(sio_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.IN(sio_in),
	.IN_H(sio_in_h),
	.TIE_LO_ESD(sio_tie_lo_esd),
	.VINREF_DFT(sio_vinref_dft),
	.VOUTREF_DFT(sio_voutref_dft),
	.DFT_REFGEN(sio_dft_refgen),
	.DM0(sio_dm0),
	.DM1(sio_dm1),
	.HLD_H_N_REFGEN(sio_hld_h_n_refgen),
	.IBUF_SEL_REFGEN(sio_ibuf_sel_refgen),
	.VOHREF(sio_vohref),
	.VOH_SEL(sio_voh_sel),
	.VREF_SEL(sio_vref_sel),
	.VREG_EN(sio_vreg_en),
	.VREG_EN_REFGEN(sio_vreg_en_refgen),
	.VTRIP_SEL_REFGEN(sio_vtrip_sel_refgen)
    );

    sky130_ef_io__gpiov2_pad gpio3_2_pad (
	.IN_H(gpio3_2_in_h),
	.IN(gpio3_2_in),
	.OUT(gpio3_2_out),
	.OE_N(gpio3_2_oe_n),
	.HLD_H_N(gpio3_2_hld_h_n),
	.ENABLE_H(gpio3_2_enable_h),
	.ENABLE_INP_H(gpio3_2_enable_inp_h),
	.ENABLE_VDDA_H(gpio3_2_enable_vdda_h),
	.ENABLE_VDDIO(gpio3_2_enable_vddio),
	.ENABLE_VSWITCH_H(gpio3_2_enable_vswitch_h),
	.INP_DIS(gpio3_2_inp_dis),
	.VTRIP_SEL(gpio3_2_vtrip_sel),
	.SLOW(gpio3_2_slow),
	.HLD_OVR(gpio3_2_hld_ovr),
	.ANALOG_EN(gpio3_2_analog_en),
	.ANALOG_SEL(gpio3_2_analog_sel),
	.ANALOG_POL(gpio3_2_analog_pol),
	.DM(gpio3_2_dm),
	.IB_MODE_SEL(gpio3_2_ib_mode_sel),
	.PAD(gpio3_2),
	.PAD_A_NOESD_H(gpio3_2_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio3_2_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio3_2_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio3_2_tie_hi_esd),
	.TIE_LO_ESD(gpio3_2_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio3_2_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio3_2_one),
	.zero(gpio3_2_zero)
    );

    sky130_ef_io__vssio_hvc_clamped_pad vssio_1_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VSSIO_PAD(vssio_1),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio5_5_pad (
	.IN_H(gpio5_5_in_h),
	.IN(gpio5_5_in),
	.OUT(gpio5_5_out),
	.OE_N(gpio5_5_oe_n),
	.HLD_H_N(gpio5_5_hld_h_n),
	.ENABLE_H(gpio5_5_enable_h),
	.ENABLE_INP_H(gpio5_5_enable_inp_h),
	.ENABLE_VDDA_H(gpio5_5_enable_vdda_h),
	.ENABLE_VDDIO(gpio5_5_enable_vddio),
	.ENABLE_VSWITCH_H(gpio5_5_enable_vswitch_h),
	.INP_DIS(gpio5_5_inp_dis),
	.VTRIP_SEL(gpio5_5_vtrip_sel),
	.SLOW(gpio5_5_slow),
	.HLD_OVR(gpio5_5_hld_ovr),
	.ANALOG_EN(gpio5_5_analog_en),
	.ANALOG_SEL(gpio5_5_analog_sel),
	.ANALOG_POL(gpio5_5_analog_pol),
	.DM(gpio5_5_dm),
	.IB_MODE_SEL(gpio5_5_ib_mode_sel),
	.PAD(gpio5_5),
	.PAD_A_NOESD_H(gpio5_5_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio5_5_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio5_5_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio5_5_tie_hi_esd),
	.TIE_LO_ESD(gpio5_5_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio5_5_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio5_5_one),
	.zero(gpio5_5_zero)
    );

    sky130_ef_io__vssd_lvc_clamped3_pad vssd1_2_pad (
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VSSD_PAD(vssd1_2),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio),
	.VCCD1(vccd1[4]),
	.VSSD1(vssd1[4])
    );

    sky130_ef_io__vssa_hvc_clamped_pad vssa3_0_pad (
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VSSA_PAD(vssa3_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__vddio_hvc_clamped_pad vddio_2_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VDDIO_PAD(vddio_2),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio2_2_pad (
	.IN_H(gpio2_2_in_h),
	.IN(gpio2_2_in),
	.OUT(gpio2_2_out),
	.OE_N(gpio2_2_oe_n),
	.HLD_H_N(gpio2_2_hld_h_n),
	.ENABLE_H(gpio2_2_enable_h),
	.ENABLE_INP_H(gpio2_2_enable_inp_h),
	.ENABLE_VDDA_H(gpio2_2_enable_vdda_h),
	.ENABLE_VDDIO(gpio2_2_enable_vddio),
	.ENABLE_VSWITCH_H(gpio2_2_enable_vswitch_h),
	.INP_DIS(gpio2_2_inp_dis),
	.VTRIP_SEL(gpio2_2_vtrip_sel),
	.SLOW(gpio2_2_slow),
	.HLD_OVR(gpio2_2_hld_ovr),
	.ANALOG_EN(gpio2_2_analog_en),
	.ANALOG_SEL(gpio2_2_analog_sel),
	.ANALOG_POL(gpio2_2_analog_pol),
	.DM(gpio2_2_dm),
	.IB_MODE_SEL(gpio2_2_ib_mode_sel),
	.PAD(gpio2_2),
	.PAD_A_NOESD_H(gpio2_2_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio2_2_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio2_2_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio2_2_tie_hi_esd),
	.TIE_LO_ESD(gpio2_2_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio2_2_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio2_2_one),
	.zero(gpio2_2_zero)
    );

    sky130_ef_io__gpiov2_pad gpio4_5_pad (
	.IN_H(gpio4_5_in_h),
	.IN(gpio4_5_in),
	.OUT(gpio4_5_out),
	.OE_N(gpio4_5_oe_n),
	.HLD_H_N(gpio4_5_hld_h_n),
	.ENABLE_H(gpio4_5_enable_h),
	.ENABLE_INP_H(gpio4_5_enable_inp_h),
	.ENABLE_VDDA_H(gpio4_5_enable_vdda_h),
	.ENABLE_VDDIO(gpio4_5_enable_vddio),
	.ENABLE_VSWITCH_H(gpio4_5_enable_vswitch_h),
	.INP_DIS(gpio4_5_inp_dis),
	.VTRIP_SEL(gpio4_5_vtrip_sel),
	.SLOW(gpio4_5_slow),
	.HLD_OVR(gpio4_5_hld_ovr),
	.ANALOG_EN(gpio4_5_analog_en),
	.ANALOG_SEL(gpio4_5_analog_sel),
	.ANALOG_POL(gpio4_5_analog_pol),
	.DM(gpio4_5_dm),
	.IB_MODE_SEL(gpio4_5_ib_mode_sel),
	.PAD(gpio4_5),
	.PAD_A_NOESD_H(gpio4_5_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio4_5_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio4_5_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio4_5_tie_hi_esd),
	.TIE_LO_ESD(gpio4_5_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio4_5_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio4_5_one),
	.zero(gpio4_5_zero)
    );

    sky130_fd_io__top_vrefcapv2 vcap_e (
	.amuxbus_a(amuxbus_a_e),
	.amuxbus_b(amuxbus_b_e),
	.cneg(vssio_q),
	.cpos(vref_e_vinref),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda1),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa1),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio)
    );

    sky130_ef_io__vssa_hvc_clamped_pad vssa2_0_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VSSA_PAD(vssa2_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__vdda_hvc_clamped_pad vdda2_1_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VDDA_PAD(vdda2_1),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_fd_io__top_gpio_ovtv2 gpio1_2_pad (
	.OUT(gpio1_2_out),
	.OE_N(gpio1_2_oe_n),
	.HLD_H_N(gpio1_2_hld_h_n),
	.ENABLE_H(gpio1_2_enable_h),
	.ENABLE_INP_H(gpio1_2_enable_inp_h),
	.ENABLE_VDDA_H(gpio1_2_enable_vdda_h),
	.ENABLE_VDDIO(gpio1_2_enable_vddio),
	.ENABLE_VSWITCH_H(gpio1_2_enable_vswitch_h),
	.INP_DIS(gpio1_2_inp_dis),
	.VTRIP_SEL(gpio1_2_vtrip_sel),
	.HYS_TRIM(gpio1_2_hys_trim),
	.SLOW(gpio1_2_slow),
	.SLEW_CTL(gpio1_2_slew_ctl),
	.HLD_OVR(gpio1_2_hld_ovr),
	.ANALOG_EN(gpio1_2_analog_en),
	.ANALOG_SEL(gpio1_2_analog_sel),
	.ANALOG_POL(gpio1_2_analog_pol),
	.DM(gpio1_2_dm),
	.IB_MODE_SEL(gpio1_2_ib_mode_sel),
	.VINREF(vref_e_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda1),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio1_2),
	.PAD_A_NOESD_H(gpio1_2_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio1_2_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio1_2_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.IN(gpio1_2_in),
	.IN_H(gpio1_2_in_h),
	.TIE_HI_ESD(gpio1_2_tie_hi_esd),
	.TIE_LO_ESD(gpio1_2_tie_lo_esd)
    );

    constant_block gpio1_2_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio1_2_one),
	.zero(gpio1_2_zero)
    );

    sky130_ef_io__gpiov2_pad gpio3_5_pad (
	.IN_H(gpio3_5_in_h),
	.IN(gpio3_5_in),
	.OUT(gpio3_5_out),
	.OE_N(gpio3_5_oe_n),
	.HLD_H_N(gpio3_5_hld_h_n),
	.ENABLE_H(gpio3_5_enable_h),
	.ENABLE_INP_H(gpio3_5_enable_inp_h),
	.ENABLE_VDDA_H(gpio3_5_enable_vdda_h),
	.ENABLE_VDDIO(gpio3_5_enable_vddio),
	.ENABLE_VSWITCH_H(gpio3_5_enable_vswitch_h),
	.INP_DIS(gpio3_5_inp_dis),
	.VTRIP_SEL(gpio3_5_vtrip_sel),
	.SLOW(gpio3_5_slow),
	.HLD_OVR(gpio3_5_hld_ovr),
	.ANALOG_EN(gpio3_5_analog_en),
	.ANALOG_SEL(gpio3_5_analog_sel),
	.ANALOG_POL(gpio3_5_analog_pol),
	.DM(gpio3_5_dm),
	.IB_MODE_SEL(gpio3_5_ib_mode_sel),
	.PAD(gpio3_5),
	.PAD_A_NOESD_H(gpio3_5_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio3_5_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio3_5_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio3_5_tie_hi_esd),
	.TIE_LO_ESD(gpio3_5_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio3_5_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio3_5_one),
	.zero(gpio3_5_zero)
    );

    sky130_ef_io__vssio_hvc_clamped_pad vssio_4_pad (
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VSSIO_PAD(vssio_4),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__vssa_hvc_clamped_pad vssa1_0_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VSSA_PAD(vssa1_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__vddio_hvc_clamped_pad vddio_5_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VDDIO_PAD(vddio_5),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__vdda_hvc_clamped_pad vdda1_1_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VDDA_PAD(vdda1_1),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio0_2_pad (
	.IN_H(gpio0_2_in_h),
	.IN(gpio0_2_in),
	.OUT(gpio0_2_out),
	.OE_N(gpio0_2_oe_n),
	.HLD_H_N(gpio0_2_hld_h_n),
	.ENABLE_H(gpio0_2_enable_h),
	.ENABLE_INP_H(gpio0_2_enable_inp_h),
	.ENABLE_VDDA_H(gpio0_2_enable_vdda_h),
	.ENABLE_VDDIO(gpio0_2_enable_vddio),
	.ENABLE_VSWITCH_H(gpio0_2_enable_vswitch_h),
	.INP_DIS(gpio0_2_inp_dis),
	.VTRIP_SEL(gpio0_2_vtrip_sel),
	.SLOW(gpio0_2_slow),
	.HLD_OVR(gpio0_2_hld_ovr),
	.ANALOG_EN(gpio0_2_analog_en),
	.ANALOG_SEL(gpio0_2_analog_sel),
	.ANALOG_POL(gpio0_2_analog_pol),
	.DM(gpio0_2_dm),
	.IB_MODE_SEL(gpio0_2_ib_mode_sel),
	.PAD(gpio0_2),
	.PAD_A_NOESD_H(gpio0_2_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio0_2_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio0_2_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio0_2_tie_hi_esd),
	.TIE_LO_ESD(gpio0_2_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio0_2_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio0_2_one),
	.zero(gpio0_2_zero)
    );

    sky130_ef_io__gpiov2_pad gpio2_5_pad (
	.IN_H(gpio2_5_in_h),
	.IN(gpio2_5_in),
	.OUT(gpio2_5_out),
	.OE_N(gpio2_5_oe_n),
	.HLD_H_N(gpio2_5_hld_h_n),
	.ENABLE_H(gpio2_5_enable_h),
	.ENABLE_INP_H(gpio2_5_enable_inp_h),
	.ENABLE_VDDA_H(gpio2_5_enable_vdda_h),
	.ENABLE_VDDIO(gpio2_5_enable_vddio),
	.ENABLE_VSWITCH_H(gpio2_5_enable_vswitch_h),
	.INP_DIS(gpio2_5_inp_dis),
	.VTRIP_SEL(gpio2_5_vtrip_sel),
	.SLOW(gpio2_5_slow),
	.HLD_OVR(gpio2_5_hld_ovr),
	.ANALOG_EN(gpio2_5_analog_en),
	.ANALOG_SEL(gpio2_5_analog_sel),
	.ANALOG_POL(gpio2_5_analog_pol),
	.DM(gpio2_5_dm),
	.IB_MODE_SEL(gpio2_5_ib_mode_sel),
	.PAD(gpio2_5),
	.PAD_A_NOESD_H(gpio2_5_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio2_5_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio2_5_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio2_5_tie_hi_esd),
	.TIE_LO_ESD(gpio2_5_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio2_5_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio2_5_one),
	.zero(gpio2_5_zero)
    );

    sky130_ef_io__vssa_hvc_clamped_pad vssa0_0_pad (
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VSSA_PAD(vssa0_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio8_1_pad (
	.IN_H(gpio8_1_in_h),
	.IN(gpio8_1_in),
	.OUT(gpio8_1_out),
	.OE_N(gpio8_1_oe_n),
	.HLD_H_N(gpio8_1_hld_h_n),
	.ENABLE_H(gpio8_1_enable_h),
	.ENABLE_INP_H(gpio8_1_enable_inp_h),
	.ENABLE_VDDA_H(gpio8_1_enable_vdda_h),
	.ENABLE_VDDIO(gpio8_1_enable_vddio),
	.ENABLE_VSWITCH_H(gpio8_1_enable_vswitch_h),
	.INP_DIS(gpio8_1_inp_dis),
	.VTRIP_SEL(gpio8_1_vtrip_sel),
	.SLOW(gpio8_1_slow),
	.HLD_OVR(gpio8_1_hld_ovr),
	.ANALOG_EN(gpio8_1_analog_en),
	.ANALOG_SEL(gpio8_1_analog_sel),
	.ANALOG_POL(gpio8_1_analog_pol),
	.DM(gpio8_1_dm),
	.IB_MODE_SEL(gpio8_1_ib_mode_sel),
	.PAD(gpio8_1),
	.PAD_A_NOESD_H(gpio8_1_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio8_1_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio8_1_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio8_1_tie_hi_esd),
	.TIE_LO_ESD(gpio8_1_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio8_1_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio8_1_one),
	.zero(gpio8_1_zero)
    );

    sky130_fd_io__top_gpio_ovtv2 gpio1_5_pad (
	.OUT(gpio1_5_out),
	.OE_N(gpio1_5_oe_n),
	.HLD_H_N(gpio1_5_hld_h_n),
	.ENABLE_H(gpio1_5_enable_h),
	.ENABLE_INP_H(gpio1_5_enable_inp_h),
	.ENABLE_VDDA_H(gpio1_5_enable_vdda_h),
	.ENABLE_VDDIO(gpio1_5_enable_vddio),
	.ENABLE_VSWITCH_H(gpio1_5_enable_vswitch_h),
	.INP_DIS(gpio1_5_inp_dis),
	.VTRIP_SEL(gpio1_5_vtrip_sel),
	.HYS_TRIM(gpio1_5_hys_trim),
	.SLOW(gpio1_5_slow),
	.SLEW_CTL(gpio1_5_slew_ctl),
	.HLD_OVR(gpio1_5_hld_ovr),
	.ANALOG_EN(gpio1_5_analog_en),
	.ANALOG_SEL(gpio1_5_analog_sel),
	.ANALOG_POL(gpio1_5_analog_pol),
	.DM(gpio1_5_dm),
	.IB_MODE_SEL(gpio1_5_ib_mode_sel),
	.VINREF(vref_e_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda1),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio1_5),
	.PAD_A_NOESD_H(gpio1_5_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio1_5_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio1_5_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.IN(gpio1_5_in),
	.IN_H(gpio1_5_in_h),
	.TIE_HI_ESD(gpio1_5_tie_hi_esd),
	.TIE_LO_ESD(gpio1_5_tie_lo_esd)
    );

    constant_block gpio1_5_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio1_5_one),
	.zero(gpio1_5_zero)
    );

    sky130_ef_io__vccd_lvc_clamped3_pad vccd2_1_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD_PAD(vccd2_1),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio),
	.VCCD1(vccd2[3]),
	.VSSD1(vssd2[3])
    );

    sky130_ef_io__vssio_hvc_clamped_pad vssio_7_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VSSIO_PAD(vssio_7),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio7_1_pad (
	.IN_H(gpio7_1_in_h),
	.IN(gpio7_1_in),
	.OUT(gpio7_1_out),
	.OE_N(gpio7_1_oe_n),
	.HLD_H_N(gpio7_1_hld_h_n),
	.ENABLE_H(gpio7_1_enable_h),
	.ENABLE_INP_H(gpio7_1_enable_inp_h),
	.ENABLE_VDDA_H(gpio7_1_enable_vdda_h),
	.ENABLE_VDDIO(gpio7_1_enable_vddio),
	.ENABLE_VSWITCH_H(gpio7_1_enable_vswitch_h),
	.INP_DIS(gpio7_1_inp_dis),
	.VTRIP_SEL(gpio7_1_vtrip_sel),
	.SLOW(gpio7_1_slow),
	.HLD_OVR(gpio7_1_hld_ovr),
	.ANALOG_EN(gpio7_1_analog_en),
	.ANALOG_SEL(gpio7_1_analog_sel),
	.ANALOG_POL(gpio7_1_analog_pol),
	.DM(gpio7_1_dm),
	.IB_MODE_SEL(gpio7_1_ib_mode_sel),
	.PAD(gpio7_1),
	.PAD_A_NOESD_H(gpio7_1_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio7_1_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio7_1_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio7_1_tie_hi_esd),
	.TIE_LO_ESD(gpio7_1_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio7_1_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio7_1_one),
	.zero(gpio7_1_zero)
    );

    sky130_ef_io__vddio_hvc_clamped_pad vddio_8_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VDDIO_PAD(vddio_8),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_fd_io__top_xres4v2 resetb_pad (
	.XRES_H_N(resetb_xres_h_n),
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.PAD(resetb),
	.PAD_A_ESD_H(resetb_pad_a_esd_h),
	.DISABLE_PULLUP_H(resetb_disable_pullup_h),
	.ENABLE_H(resetb_enable_h),
	.EN_VDDIO_SIG_H(resetb_en_vddio_sig_h),
	.INP_SEL_H(resetb_inp_sel_h),
	.FILT_IN_H(resetb_filt_in_h),
	.PULLUP_H(resetb_pullup_h),
	.ENABLE_VDDIO(resetb_enable_vddio),
	.TIE_LO_ESD(resetb_tie_lo_esd),
	.TIE_HI_ESD(resetb_tie_hi_esd),
	.TIE_WEAK_HI_H(resetb_tie_weak_hi_h),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio0_5_pad (
	.IN_H(gpio0_5_in_h),
	.IN(gpio0_5_in),
	.OUT(gpio0_5_out),
	.OE_N(gpio0_5_oe_n),
	.HLD_H_N(gpio0_5_hld_h_n),
	.ENABLE_H(gpio0_5_enable_h),
	.ENABLE_INP_H(gpio0_5_enable_inp_h),
	.ENABLE_VDDA_H(gpio0_5_enable_vdda_h),
	.ENABLE_VDDIO(gpio0_5_enable_vddio),
	.ENABLE_VSWITCH_H(gpio0_5_enable_vswitch_h),
	.INP_DIS(gpio0_5_inp_dis),
	.VTRIP_SEL(gpio0_5_vtrip_sel),
	.SLOW(gpio0_5_slow),
	.HLD_OVR(gpio0_5_hld_ovr),
	.ANALOG_EN(gpio0_5_analog_en),
	.ANALOG_SEL(gpio0_5_analog_sel),
	.ANALOG_POL(gpio0_5_analog_pol),
	.DM(gpio0_5_dm),
	.IB_MODE_SEL(gpio0_5_ib_mode_sel),
	.PAD(gpio0_5),
	.PAD_A_NOESD_H(gpio0_5_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio0_5_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio0_5_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio0_5_tie_hi_esd),
	.TIE_LO_ESD(gpio0_5_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio0_5_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio0_5_one),
	.zero(gpio0_5_zero)
    );

    sky130_ef_io__vccd_lvc_clamped3_pad vccd1_1_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD_PAD(vccd1_1),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio),
	.VCCD1(vccd1[3]),
	.VSSD1(vssd1[3])
    );

    sky130_fd_io__top_gpio_ovtv2 gpio6_1_pad (
	.OUT(gpio6_1_out),
	.OE_N(gpio6_1_oe_n),
	.HLD_H_N(gpio6_1_hld_h_n),
	.ENABLE_H(gpio6_1_enable_h),
	.ENABLE_INP_H(gpio6_1_enable_inp_h),
	.ENABLE_VDDA_H(gpio6_1_enable_vdda_h),
	.ENABLE_VDDIO(gpio6_1_enable_vddio),
	.ENABLE_VSWITCH_H(gpio6_1_enable_vswitch_h),
	.INP_DIS(gpio6_1_inp_dis),
	.VTRIP_SEL(gpio6_1_vtrip_sel),
	.HYS_TRIM(gpio6_1_hys_trim),
	.SLOW(gpio6_1_slow),
	.SLEW_CTL(gpio6_1_slew_ctl),
	.HLD_OVR(gpio6_1_hld_ovr),
	.ANALOG_EN(gpio6_1_analog_en),
	.ANALOG_SEL(gpio6_1_analog_sel),
	.ANALOG_POL(gpio6_1_analog_pol),
	.DM(gpio6_1_dm),
	.IB_MODE_SEL(gpio6_1_ib_mode_sel),
	.VINREF(vref_w_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda2),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio6_1),
	.PAD_A_NOESD_H(gpio6_1_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio6_1_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio6_1_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.IN(gpio6_1_in),
	.IN_H(gpio6_1_in_h),
	.TIE_HI_ESD(gpio6_1_tie_hi_esd),
	.TIE_LO_ESD(gpio6_1_tie_lo_esd)
    );

    constant_block gpio6_1_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio6_1_one),
	.zero(gpio6_1_zero)
    );

    sky130_ef_io__gpiov2_pad gpio8_4_pad (
	.IN_H(gpio8_4_in_h),
	.IN(gpio8_4_in),
	.OUT(gpio8_4_out),
	.OE_N(gpio8_4_oe_n),
	.HLD_H_N(gpio8_4_hld_h_n),
	.ENABLE_H(gpio8_4_enable_h),
	.ENABLE_INP_H(gpio8_4_enable_inp_h),
	.ENABLE_VDDA_H(gpio8_4_enable_vdda_h),
	.ENABLE_VDDIO(gpio8_4_enable_vddio),
	.ENABLE_VSWITCH_H(gpio8_4_enable_vswitch_h),
	.INP_DIS(gpio8_4_inp_dis),
	.VTRIP_SEL(gpio8_4_vtrip_sel),
	.SLOW(gpio8_4_slow),
	.HLD_OVR(gpio8_4_hld_ovr),
	.ANALOG_EN(gpio8_4_analog_en),
	.ANALOG_SEL(gpio8_4_analog_sel),
	.ANALOG_POL(gpio8_4_analog_pol),
	.DM(gpio8_4_dm),
	.IB_MODE_SEL(gpio8_4_ib_mode_sel),
	.PAD(gpio8_4),
	.PAD_A_NOESD_H(gpio8_4_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio8_4_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio8_4_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio8_4_tie_hi_esd),
	.TIE_LO_ESD(gpio8_4_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio8_4_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio8_4_one),
	.zero(gpio8_4_zero)
    );

    sky130_ef_io__vccd_lvc_clamped_pad vccd0_1_pad (
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VCCD_PAD(vccd0_1),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio5_1_pad (
	.IN_H(gpio5_1_in_h),
	.IN(gpio5_1_in),
	.OUT(gpio5_1_out),
	.OE_N(gpio5_1_oe_n),
	.HLD_H_N(gpio5_1_hld_h_n),
	.ENABLE_H(gpio5_1_enable_h),
	.ENABLE_INP_H(gpio5_1_enable_inp_h),
	.ENABLE_VDDA_H(gpio5_1_enable_vdda_h),
	.ENABLE_VDDIO(gpio5_1_enable_vddio),
	.ENABLE_VSWITCH_H(gpio5_1_enable_vswitch_h),
	.INP_DIS(gpio5_1_inp_dis),
	.VTRIP_SEL(gpio5_1_vtrip_sel),
	.SLOW(gpio5_1_slow),
	.HLD_OVR(gpio5_1_hld_ovr),
	.ANALOG_EN(gpio5_1_analog_en),
	.ANALOG_SEL(gpio5_1_analog_sel),
	.ANALOG_POL(gpio5_1_analog_pol),
	.DM(gpio5_1_dm),
	.IB_MODE_SEL(gpio5_1_ib_mode_sel),
	.PAD(gpio5_1),
	.PAD_A_NOESD_H(gpio5_1_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio5_1_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio5_1_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio5_1_tie_hi_esd),
	.TIE_LO_ESD(gpio5_1_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio5_1_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio5_1_one),
	.zero(gpio5_1_zero)
    );

    sky130_ef_io__gpiov2_pad gpio7_4_pad (
	.IN_H(gpio7_4_in_h),
	.IN(gpio7_4_in),
	.OUT(gpio7_4_out),
	.OE_N(gpio7_4_oe_n),
	.HLD_H_N(gpio7_4_hld_h_n),
	.ENABLE_H(gpio7_4_enable_h),
	.ENABLE_INP_H(gpio7_4_enable_inp_h),
	.ENABLE_VDDA_H(gpio7_4_enable_vdda_h),
	.ENABLE_VDDIO(gpio7_4_enable_vddio),
	.ENABLE_VSWITCH_H(gpio7_4_enable_vswitch_h),
	.INP_DIS(gpio7_4_inp_dis),
	.VTRIP_SEL(gpio7_4_vtrip_sel),
	.SLOW(gpio7_4_slow),
	.HLD_OVR(gpio7_4_hld_ovr),
	.ANALOG_EN(gpio7_4_analog_en),
	.ANALOG_SEL(gpio7_4_analog_sel),
	.ANALOG_POL(gpio7_4_analog_pol),
	.DM(gpio7_4_dm),
	.IB_MODE_SEL(gpio7_4_ib_mode_sel),
	.PAD(gpio7_4),
	.PAD_A_NOESD_H(gpio7_4_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio7_4_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio7_4_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio7_4_tie_hi_esd),
	.TIE_LO_ESD(gpio7_4_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio7_4_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio7_4_one),
	.zero(gpio7_4_zero)
    );

    sky130_fd_io__top_gpiovrefv2 vref_e (
	.amuxbus_a(amuxbus_a_e),
	.amuxbus_b(amuxbus_b_e),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda1),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa1),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio),
	.enable_h(vref_e_enable_h),
	.hld_h_n(vref_e_hld_h_n),
	.ref_sel(vref_e_ref_sel),
	.vrefgen_en(vref_e_vrefgen_en),
	.vinref(vref_e_vinref)
    );

    sky130_fd_io__top_amuxsplitv2 muxsplit_sw (
	.amuxbus_a_l(amuxbus_a_s),
	.amuxbus_a_r(amuxbus_a_w),
	.amuxbus_b_l(amuxbus_b_s),
	.amuxbus_b_r(amuxbus_b_w),
	.enable_vdda_h(muxsplit_sw_enable_vdda_h),
	.hld_vdda_h_n(muxsplit_sw_hld_vdda_h_n),
	.switch_aa_s0(muxsplit_sw_switch_aa_s0),
	.switch_aa_sl(muxsplit_sw_switch_aa_sl),
	.switch_aa_sr(muxsplit_sw_switch_aa_sr),
	.switch_bb_s0(muxsplit_sw_switch_bb_s0),
	.switch_bb_sl(muxsplit_sw_switch_bb_sl),
	.switch_bb_sr(muxsplit_sw_switch_bb_sr),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda3),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa3),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio4_1_pad (
	.IN_H(gpio4_1_in_h),
	.IN(gpio4_1_in),
	.OUT(gpio4_1_out),
	.OE_N(gpio4_1_oe_n),
	.HLD_H_N(gpio4_1_hld_h_n),
	.ENABLE_H(gpio4_1_enable_h),
	.ENABLE_INP_H(gpio4_1_enable_inp_h),
	.ENABLE_VDDA_H(gpio4_1_enable_vdda_h),
	.ENABLE_VDDIO(gpio4_1_enable_vddio),
	.ENABLE_VSWITCH_H(gpio4_1_enable_vswitch_h),
	.INP_DIS(gpio4_1_inp_dis),
	.VTRIP_SEL(gpio4_1_vtrip_sel),
	.SLOW(gpio4_1_slow),
	.HLD_OVR(gpio4_1_hld_ovr),
	.ANALOG_EN(gpio4_1_analog_en),
	.ANALOG_SEL(gpio4_1_analog_sel),
	.ANALOG_POL(gpio4_1_analog_pol),
	.DM(gpio4_1_dm),
	.IB_MODE_SEL(gpio4_1_ib_mode_sel),
	.PAD(gpio4_1),
	.PAD_A_NOESD_H(gpio4_1_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio4_1_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio4_1_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio4_1_tie_hi_esd),
	.TIE_LO_ESD(gpio4_1_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio4_1_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio4_1_one),
	.zero(gpio4_1_zero)
    );

    sky130_ef_io__vssd_lvc_clamped3_pad vssd2_1_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VSSD_PAD(vssd2_1),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio),
	.VCCD1(vccd2[2]),
	.VSSD1(vssd2[2])
    );

    sky130_fd_io__top_gpio_ovtv2 gpio6_4_pad (
	.OUT(gpio6_4_out),
	.OE_N(gpio6_4_oe_n),
	.HLD_H_N(gpio6_4_hld_h_n),
	.ENABLE_H(gpio6_4_enable_h),
	.ENABLE_INP_H(gpio6_4_enable_inp_h),
	.ENABLE_VDDA_H(gpio6_4_enable_vdda_h),
	.ENABLE_VDDIO(gpio6_4_enable_vddio),
	.ENABLE_VSWITCH_H(gpio6_4_enable_vswitch_h),
	.INP_DIS(gpio6_4_inp_dis),
	.VTRIP_SEL(gpio6_4_vtrip_sel),
	.HYS_TRIM(gpio6_4_hys_trim),
	.SLOW(gpio6_4_slow),
	.SLEW_CTL(gpio6_4_slew_ctl),
	.HLD_OVR(gpio6_4_hld_ovr),
	.ANALOG_EN(gpio6_4_analog_en),
	.ANALOG_SEL(gpio6_4_analog_sel),
	.ANALOG_POL(gpio6_4_analog_pol),
	.DM(gpio6_4_dm),
	.IB_MODE_SEL(gpio6_4_ib_mode_sel),
	.VINREF(vref_w_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda2),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio6_4),
	.PAD_A_NOESD_H(gpio6_4_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio6_4_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio6_4_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.IN(gpio6_4_in),
	.IN_H(gpio6_4_in_h),
	.TIE_HI_ESD(gpio6_4_tie_hi_esd),
	.TIE_LO_ESD(gpio6_4_tie_lo_esd)
    );

    constant_block gpio6_4_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio6_4_one),
	.zero(gpio6_4_zero)
    );

    sky130_ef_io__gpiov2_pad gpio8_7_pad (
	.IN_H(gpio8_7_in_h),
	.IN(gpio8_7_in),
	.OUT(gpio8_7_out),
	.OE_N(gpio8_7_oe_n),
	.HLD_H_N(gpio8_7_hld_h_n),
	.ENABLE_H(gpio8_7_enable_h),
	.ENABLE_INP_H(gpio8_7_enable_inp_h),
	.ENABLE_VDDA_H(gpio8_7_enable_vdda_h),
	.ENABLE_VDDIO(gpio8_7_enable_vddio),
	.ENABLE_VSWITCH_H(gpio8_7_enable_vswitch_h),
	.INP_DIS(gpio8_7_inp_dis),
	.VTRIP_SEL(gpio8_7_vtrip_sel),
	.SLOW(gpio8_7_slow),
	.HLD_OVR(gpio8_7_hld_ovr),
	.ANALOG_EN(gpio8_7_analog_en),
	.ANALOG_SEL(gpio8_7_analog_sel),
	.ANALOG_POL(gpio8_7_analog_pol),
	.DM(gpio8_7_dm),
	.IB_MODE_SEL(gpio8_7_ib_mode_sel),
	.PAD(gpio8_7),
	.PAD_A_NOESD_H(gpio8_7_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio8_7_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio8_7_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio8_7_tie_hi_esd),
	.TIE_LO_ESD(gpio8_7_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio8_7_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio8_7_one),
	.zero(gpio8_7_zero)
    );

    sky130_fd_io__top_pwrdetv2 pwrdet_s (
	.out1_vddd_hv(pwrdet_out1_vddd_hv),
	.out1_vddio_hv(pwrdet_out1_vddio_hv),
	.out2_vddd_hv(pwrdet_out2_vddd_hv),
	.out2_vddio_hv(pwrdet_out2_vddio_hv),
	.out3_vddd_hv(pwrdet_out3_vddd_hv),
	.out3_vddio_hv(pwrdet_out3_vddio_hv),
	.tie_lo_esd(pwrdet_tie_lo_esd),
	.vddd_present_vddio_hv(pwrdet_vddd_present_vddio_hv),
	.vddio_present_vddd_hv(pwrdet_vddio_present_vddd_hv),
	.in1_vddd_hv(pwrdet_in1_vddd_hv),
	.in1_vddio_hv(pwrdet_in1_vddio_hv),
	.in2_vddd_hv(pwrdet_in2_vddd_hv),
	.in2_vddio_hv(pwrdet_in2_vddio_hv),
	.in3_vddd_hv(pwrdet_in3_vddd_hv),
	.in3_vddio_hv(pwrdet_in3_vddio_hv),
	.rst_por_hv_n(pwrdet_rst_por_hv_n),
	.vccd(vccd0),
	.vddd1(vdda3),
	.vddd2(vdda3),
	.vssa(vssa3),
	.vssd(vssd0),
	.vddio_q(vddio_q),
	.vssio_q()		// This pin has no physical connection.
    );

    sky130_ef_io__gpiov2_pad gpio3_1_pad (
	.IN_H(gpio3_1_in_h),
	.IN(gpio3_1_in),
	.OUT(gpio3_1_out),
	.OE_N(gpio3_1_oe_n),
	.HLD_H_N(gpio3_1_hld_h_n),
	.ENABLE_H(gpio3_1_enable_h),
	.ENABLE_INP_H(gpio3_1_enable_inp_h),
	.ENABLE_VDDA_H(gpio3_1_enable_vdda_h),
	.ENABLE_VDDIO(gpio3_1_enable_vddio),
	.ENABLE_VSWITCH_H(gpio3_1_enable_vswitch_h),
	.INP_DIS(gpio3_1_inp_dis),
	.VTRIP_SEL(gpio3_1_vtrip_sel),
	.SLOW(gpio3_1_slow),
	.HLD_OVR(gpio3_1_hld_ovr),
	.ANALOG_EN(gpio3_1_analog_en),
	.ANALOG_SEL(gpio3_1_analog_sel),
	.ANALOG_POL(gpio3_1_analog_pol),
	.DM(gpio3_1_dm),
	.IB_MODE_SEL(gpio3_1_ib_mode_sel),
	.PAD(gpio3_1),
	.PAD_A_NOESD_H(gpio3_1_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio3_1_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio3_1_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio3_1_tie_hi_esd),
	.TIE_LO_ESD(gpio3_1_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio3_1_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio3_1_one),
	.zero(gpio3_1_zero)
    );

    sky130_ef_io__vssio_hvc_clamped_pad vssio_0_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VSSIO_PAD(vssio_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio5_4_pad (
	.IN_H(gpio5_4_in_h),
	.IN(gpio5_4_in),
	.OUT(gpio5_4_out),
	.OE_N(gpio5_4_oe_n),
	.HLD_H_N(gpio5_4_hld_h_n),
	.ENABLE_H(gpio5_4_enable_h),
	.ENABLE_INP_H(gpio5_4_enable_inp_h),
	.ENABLE_VDDA_H(gpio5_4_enable_vdda_h),
	.ENABLE_VDDIO(gpio5_4_enable_vddio),
	.ENABLE_VSWITCH_H(gpio5_4_enable_vswitch_h),
	.INP_DIS(gpio5_4_inp_dis),
	.VTRIP_SEL(gpio5_4_vtrip_sel),
	.SLOW(gpio5_4_slow),
	.HLD_OVR(gpio5_4_hld_ovr),
	.ANALOG_EN(gpio5_4_analog_en),
	.ANALOG_SEL(gpio5_4_analog_sel),
	.ANALOG_POL(gpio5_4_analog_pol),
	.DM(gpio5_4_dm),
	.IB_MODE_SEL(gpio5_4_ib_mode_sel),
	.PAD(gpio5_4),
	.PAD_A_NOESD_H(gpio5_4_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio5_4_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio5_4_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio5_4_tie_hi_esd),
	.TIE_LO_ESD(gpio5_4_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio5_4_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio5_4_one),
	.zero(gpio5_4_zero)
    );

    sky130_ef_io__vssd_lvc_clamped3_pad vssd1_1_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VSSD_PAD(vssd1_1),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio),
	.VCCD1(vccd1[2]),
	.VSSD1(vssd1[2])
    );

    sky130_ef_io__gpiov2_pad gpio7_7_pad (
	.IN_H(gpio7_7_in_h),
	.IN(gpio7_7_in),
	.OUT(gpio7_7_out),
	.OE_N(gpio7_7_oe_n),
	.HLD_H_N(gpio7_7_hld_h_n),
	.ENABLE_H(gpio7_7_enable_h),
	.ENABLE_INP_H(gpio7_7_enable_inp_h),
	.ENABLE_VDDA_H(gpio7_7_enable_vdda_h),
	.ENABLE_VDDIO(gpio7_7_enable_vddio),
	.ENABLE_VSWITCH_H(gpio7_7_enable_vswitch_h),
	.INP_DIS(gpio7_7_inp_dis),
	.VTRIP_SEL(gpio7_7_vtrip_sel),
	.SLOW(gpio7_7_slow),
	.HLD_OVR(gpio7_7_hld_ovr),
	.ANALOG_EN(gpio7_7_analog_en),
	.ANALOG_SEL(gpio7_7_analog_sel),
	.ANALOG_POL(gpio7_7_analog_pol),
	.DM(gpio7_7_dm),
	.IB_MODE_SEL(gpio7_7_ib_mode_sel),
	.PAD(gpio7_7),
	.PAD_A_NOESD_H(gpio7_7_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio7_7_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio7_7_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio7_7_tie_hi_esd),
	.TIE_LO_ESD(gpio7_7_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio7_7_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio7_7_one),
	.zero(gpio7_7_zero)
    );

    sky130_ef_io__vddio_hvc_clamped_pad vddio_1_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VDDIO_PAD(vddio_1),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__vdda_hvc_clamped_pad vdda3_0_pad (
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VDDA_PAD(vdda3_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio2_1_pad (
	.IN_H(gpio2_1_in_h),
	.IN(gpio2_1_in),
	.OUT(gpio2_1_out),
	.OE_N(gpio2_1_oe_n),
	.HLD_H_N(gpio2_1_hld_h_n),
	.ENABLE_H(gpio2_1_enable_h),
	.ENABLE_INP_H(gpio2_1_enable_inp_h),
	.ENABLE_VDDA_H(gpio2_1_enable_vdda_h),
	.ENABLE_VDDIO(gpio2_1_enable_vddio),
	.ENABLE_VSWITCH_H(gpio2_1_enable_vswitch_h),
	.INP_DIS(gpio2_1_inp_dis),
	.VTRIP_SEL(gpio2_1_vtrip_sel),
	.SLOW(gpio2_1_slow),
	.HLD_OVR(gpio2_1_hld_ovr),
	.ANALOG_EN(gpio2_1_analog_en),
	.ANALOG_SEL(gpio2_1_analog_sel),
	.ANALOG_POL(gpio2_1_analog_pol),
	.DM(gpio2_1_dm),
	.IB_MODE_SEL(gpio2_1_ib_mode_sel),
	.PAD(gpio2_1),
	.PAD_A_NOESD_H(gpio2_1_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio2_1_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio2_1_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio2_1_tie_hi_esd),
	.TIE_LO_ESD(gpio2_1_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio2_1_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio2_1_one),
	.zero(gpio2_1_zero)
    );

    sky130_ef_io__gpiov2_pad gpio4_4_pad (
	.IN_H(gpio4_4_in_h),
	.IN(gpio4_4_in),
	.OUT(gpio4_4_out),
	.OE_N(gpio4_4_oe_n),
	.HLD_H_N(gpio4_4_hld_h_n),
	.ENABLE_H(gpio4_4_enable_h),
	.ENABLE_INP_H(gpio4_4_enable_inp_h),
	.ENABLE_VDDA_H(gpio4_4_enable_vdda_h),
	.ENABLE_VDDIO(gpio4_4_enable_vddio),
	.ENABLE_VSWITCH_H(gpio4_4_enable_vswitch_h),
	.INP_DIS(gpio4_4_inp_dis),
	.VTRIP_SEL(gpio4_4_vtrip_sel),
	.SLOW(gpio4_4_slow),
	.HLD_OVR(gpio4_4_hld_ovr),
	.ANALOG_EN(gpio4_4_analog_en),
	.ANALOG_SEL(gpio4_4_analog_sel),
	.ANALOG_POL(gpio4_4_analog_pol),
	.DM(gpio4_4_dm),
	.IB_MODE_SEL(gpio4_4_ib_mode_sel),
	.PAD(gpio4_4),
	.PAD_A_NOESD_H(gpio4_4_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio4_4_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio4_4_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio4_4_tie_hi_esd),
	.TIE_LO_ESD(gpio4_4_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio4_4_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio4_4_one),
	.zero(gpio4_4_zero)
    );

    sky130_ef_io__vssd_lvc_clamped_pad vssd0_1_pad (
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VSSD_PAD(vssd0_1),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad select_pad (
	.IN_H(select_in_h),
	.IN(select_in),
	.OUT(select_out),
	.OE_N(select_oe_n),
	.HLD_H_N(select_hld_h_n),
	.ENABLE_H(select_enable_h),
	.ENABLE_INP_H(select_enable_inp_h),
	.ENABLE_VDDA_H(select_enable_vdda_h),
	.ENABLE_VDDIO(select_enable_vddio),
	.ENABLE_VSWITCH_H(select_enable_vswitch_h),
	.INP_DIS(select_inp_dis),
	.VTRIP_SEL(select_vtrip_sel),
	.SLOW(select_slow),
	.HLD_OVR(select_hld_ovr),
	.ANALOG_EN(select_analog_en),
	.ANALOG_SEL(select_analog_sel),
	.ANALOG_POL(select_analog_pol),
	.DM(select_dm),
	.IB_MODE_SEL(select_ib_mode_sel),
	.PAD(select),
	.PAD_A_NOESD_H(select_pad_a_noesd_h),
	.PAD_A_ESD_0_H(select_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(select_pad_a_esd_1_h),
	.TIE_HI_ESD(select_tie_hi_esd),
	.TIE_LO_ESD(select_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block select_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(select_one),
	.zero(select_zero)
    );

    sky130_fd_io__top_gpio_ovtv2 gpio6_7_pad (
	.OUT(gpio6_7_out),
	.OE_N(gpio6_7_oe_n),
	.HLD_H_N(gpio6_7_hld_h_n),
	.ENABLE_H(gpio6_7_enable_h),
	.ENABLE_INP_H(gpio6_7_enable_inp_h),
	.ENABLE_VDDA_H(gpio6_7_enable_vdda_h),
	.ENABLE_VDDIO(gpio6_7_enable_vddio),
	.ENABLE_VSWITCH_H(gpio6_7_enable_vswitch_h),
	.INP_DIS(gpio6_7_inp_dis),
	.VTRIP_SEL(gpio6_7_vtrip_sel),
	.HYS_TRIM(gpio6_7_hys_trim),
	.SLOW(gpio6_7_slow),
	.SLEW_CTL(gpio6_7_slew_ctl),
	.HLD_OVR(gpio6_7_hld_ovr),
	.ANALOG_EN(gpio6_7_analog_en),
	.ANALOG_SEL(gpio6_7_analog_sel),
	.ANALOG_POL(gpio6_7_analog_pol),
	.DM(gpio6_7_dm),
	.IB_MODE_SEL(gpio6_7_ib_mode_sel),
	.VINREF(vref_w_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda2),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio6_7),
	.PAD_A_NOESD_H(gpio6_7_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio6_7_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio6_7_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.IN(gpio6_7_in),
	.IN_H(gpio6_7_in_h),
	.TIE_HI_ESD(gpio6_7_tie_hi_esd),
	.TIE_LO_ESD(gpio6_7_tie_lo_esd)
    );

    constant_block gpio6_7_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio6_7_one),
	.zero(gpio6_7_zero)
    );

    sky130_fd_io__top_analog_pad xi1_pad (
	.pad_core(xi1_core),
	.pad(xi1),
	.amuxbus_a(amuxbus_a_s),
	.amuxbus_b(amuxbus_b_s),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda3),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa3),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio)
    );

    sky130_ef_io__vdda_hvc_clamped_pad vdda2_0_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VDDA_PAD(vdda2_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_fd_io__top_gpio_ovtv2 gpio1_1_pad (
	.OUT(gpio1_1_out),
	.OE_N(gpio1_1_oe_n),
	.HLD_H_N(gpio1_1_hld_h_n),
	.ENABLE_H(gpio1_1_enable_h),
	.ENABLE_INP_H(gpio1_1_enable_inp_h),
	.ENABLE_VDDA_H(gpio1_1_enable_vdda_h),
	.ENABLE_VDDIO(gpio1_1_enable_vddio),
	.ENABLE_VSWITCH_H(gpio1_1_enable_vswitch_h),
	.INP_DIS(gpio1_1_inp_dis),
	.VTRIP_SEL(gpio1_1_vtrip_sel),
	.HYS_TRIM(gpio1_1_hys_trim),
	.SLOW(gpio1_1_slow),
	.SLEW_CTL(gpio1_1_slew_ctl),
	.HLD_OVR(gpio1_1_hld_ovr),
	.ANALOG_EN(gpio1_1_analog_en),
	.ANALOG_SEL(gpio1_1_analog_sel),
	.ANALOG_POL(gpio1_1_analog_pol),
	.DM(gpio1_1_dm),
	.IB_MODE_SEL(gpio1_1_ib_mode_sel),
	.VINREF(vref_e_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda1),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio1_1),
	.PAD_A_NOESD_H(gpio1_1_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio1_1_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio1_1_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.IN(gpio1_1_in),
	.IN_H(gpio1_1_in_h),
	.TIE_HI_ESD(gpio1_1_tie_hi_esd),
	.TIE_LO_ESD(gpio1_1_tie_lo_esd)
    );

    constant_block gpio1_1_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio1_1_one),
	.zero(gpio1_1_zero)
    );

    sky130_ef_io__vssio_hvc_clamped_pad vssio_3_pad (
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VSSIO_PAD(vssio_3),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio3_4_pad (
	.IN_H(gpio3_4_in_h),
	.IN(gpio3_4_in),
	.OUT(gpio3_4_out),
	.OE_N(gpio3_4_oe_n),
	.HLD_H_N(gpio3_4_hld_h_n),
	.ENABLE_H(gpio3_4_enable_h),
	.ENABLE_INP_H(gpio3_4_enable_inp_h),
	.ENABLE_VDDA_H(gpio3_4_enable_vdda_h),
	.ENABLE_VDDIO(gpio3_4_enable_vddio),
	.ENABLE_VSWITCH_H(gpio3_4_enable_vswitch_h),
	.INP_DIS(gpio3_4_inp_dis),
	.VTRIP_SEL(gpio3_4_vtrip_sel),
	.SLOW(gpio3_4_slow),
	.HLD_OVR(gpio3_4_hld_ovr),
	.ANALOG_EN(gpio3_4_analog_en),
	.ANALOG_SEL(gpio3_4_analog_sel),
	.ANALOG_POL(gpio3_4_analog_pol),
	.DM(gpio3_4_dm),
	.IB_MODE_SEL(gpio3_4_ib_mode_sel),
	.PAD(gpio3_4),
	.PAD_A_NOESD_H(gpio3_4_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio3_4_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio3_4_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio3_4_tie_hi_esd),
	.TIE_LO_ESD(gpio3_4_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio3_4_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio3_4_one),
	.zero(gpio3_4_zero)
    );

    sky130_ef_io__gpiov2_pad gpio5_7_pad (
	.IN_H(gpio5_7_in_h),
	.IN(gpio5_7_in),
	.OUT(gpio5_7_out),
	.OE_N(gpio5_7_oe_n),
	.HLD_H_N(gpio5_7_hld_h_n),
	.ENABLE_H(gpio5_7_enable_h),
	.ENABLE_INP_H(gpio5_7_enable_inp_h),
	.ENABLE_VDDA_H(gpio5_7_enable_vdda_h),
	.ENABLE_VDDIO(gpio5_7_enable_vddio),
	.ENABLE_VSWITCH_H(gpio5_7_enable_vswitch_h),
	.INP_DIS(gpio5_7_inp_dis),
	.VTRIP_SEL(gpio5_7_vtrip_sel),
	.SLOW(gpio5_7_slow),
	.HLD_OVR(gpio5_7_hld_ovr),
	.ANALOG_EN(gpio5_7_analog_en),
	.ANALOG_SEL(gpio5_7_analog_sel),
	.ANALOG_POL(gpio5_7_analog_pol),
	.DM(gpio5_7_dm),
	.IB_MODE_SEL(gpio5_7_ib_mode_sel),
	.PAD(gpio5_7),
	.PAD_A_NOESD_H(gpio5_7_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio5_7_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio5_7_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio5_7_tie_hi_esd),
	.TIE_LO_ESD(gpio5_7_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio5_7_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio5_7_one),
	.zero(gpio5_7_zero)
    );

    sky130_ef_io__vddio_hvc_clamped_pad vddio_4_pad (
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VDDIO_PAD(vddio_4),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_fd_io__top_amuxsplitv2 muxsplit_nw (
	.amuxbus_a_l(amuxbus_a_w),
	.amuxbus_a_r(amuxbus_a_n),
	.amuxbus_b_l(amuxbus_b_w),
	.amuxbus_b_r(amuxbus_b_n),
	.enable_vdda_h(muxsplit_nw_enable_vdda_h),
	.hld_vdda_h_n(muxsplit_nw_hld_vdda_h_n),
	.switch_aa_s0(muxsplit_nw_switch_aa_s0),
	.switch_aa_sl(muxsplit_nw_switch_aa_sl),
	.switch_aa_sr(muxsplit_nw_switch_aa_sr),
	.switch_bb_s0(muxsplit_nw_switch_bb_s0),
	.switch_bb_sl(muxsplit_nw_switch_bb_sl),
	.switch_bb_sr(muxsplit_nw_switch_bb_sr),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda0),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa0),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio0_1_pad (
	.IN_H(gpio0_1_in_h),
	.IN(gpio0_1_in),
	.OUT(gpio0_1_out),
	.OE_N(gpio0_1_oe_n),
	.HLD_H_N(gpio0_1_hld_h_n),
	.ENABLE_H(gpio0_1_enable_h),
	.ENABLE_INP_H(gpio0_1_enable_inp_h),
	.ENABLE_VDDA_H(gpio0_1_enable_vdda_h),
	.ENABLE_VDDIO(gpio0_1_enable_vddio),
	.ENABLE_VSWITCH_H(gpio0_1_enable_vswitch_h),
	.INP_DIS(gpio0_1_inp_dis),
	.VTRIP_SEL(gpio0_1_vtrip_sel),
	.SLOW(gpio0_1_slow),
	.HLD_OVR(gpio0_1_hld_ovr),
	.ANALOG_EN(gpio0_1_analog_en),
	.ANALOG_SEL(gpio0_1_analog_sel),
	.ANALOG_POL(gpio0_1_analog_pol),
	.DM(gpio0_1_dm),
	.IB_MODE_SEL(gpio0_1_ib_mode_sel),
	.PAD(gpio0_1),
	.PAD_A_NOESD_H(gpio0_1_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio0_1_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio0_1_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio0_1_tie_hi_esd),
	.TIE_LO_ESD(gpio0_1_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio0_1_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio0_1_one),
	.zero(gpio0_1_zero)
    );

    sky130_ef_io__vdda_hvc_clamped_pad vdda1_0_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VDDA_PAD(vdda1_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio2_4_pad (
	.IN_H(gpio2_4_in_h),
	.IN(gpio2_4_in),
	.OUT(gpio2_4_out),
	.OE_N(gpio2_4_oe_n),
	.HLD_H_N(gpio2_4_hld_h_n),
	.ENABLE_H(gpio2_4_enable_h),
	.ENABLE_INP_H(gpio2_4_enable_inp_h),
	.ENABLE_VDDA_H(gpio2_4_enable_vdda_h),
	.ENABLE_VDDIO(gpio2_4_enable_vddio),
	.ENABLE_VSWITCH_H(gpio2_4_enable_vswitch_h),
	.INP_DIS(gpio2_4_inp_dis),
	.VTRIP_SEL(gpio2_4_vtrip_sel),
	.SLOW(gpio2_4_slow),
	.HLD_OVR(gpio2_4_hld_ovr),
	.ANALOG_EN(gpio2_4_analog_en),
	.ANALOG_SEL(gpio2_4_analog_sel),
	.ANALOG_POL(gpio2_4_analog_pol),
	.DM(gpio2_4_dm),
	.IB_MODE_SEL(gpio2_4_ib_mode_sel),
	.PAD(gpio2_4),
	.PAD_A_NOESD_H(gpio2_4_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio2_4_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio2_4_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio2_4_tie_hi_esd),
	.TIE_LO_ESD(gpio2_4_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio2_4_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio2_4_one),
	.zero(gpio2_4_zero)
    );

    sky130_ef_io__gpiov2_pad gpio4_7_pad (
	.IN_H(gpio4_7_in_h),
	.IN(gpio4_7_in),
	.OUT(gpio4_7_out),
	.OE_N(gpio4_7_oe_n),
	.HLD_H_N(gpio4_7_hld_h_n),
	.ENABLE_H(gpio4_7_enable_h),
	.ENABLE_INP_H(gpio4_7_enable_inp_h),
	.ENABLE_VDDA_H(gpio4_7_enable_vdda_h),
	.ENABLE_VDDIO(gpio4_7_enable_vddio),
	.ENABLE_VSWITCH_H(gpio4_7_enable_vswitch_h),
	.INP_DIS(gpio4_7_inp_dis),
	.VTRIP_SEL(gpio4_7_vtrip_sel),
	.SLOW(gpio4_7_slow),
	.HLD_OVR(gpio4_7_hld_ovr),
	.ANALOG_EN(gpio4_7_analog_en),
	.ANALOG_SEL(gpio4_7_analog_sel),
	.ANALOG_POL(gpio4_7_analog_pol),
	.DM(gpio4_7_dm),
	.IB_MODE_SEL(gpio4_7_ib_mode_sel),
	.PAD(gpio4_7),
	.PAD_A_NOESD_H(gpio4_7_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio4_7_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio4_7_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio4_7_tie_hi_esd),
	.TIE_LO_ESD(gpio4_7_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio4_7_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio4_7_one),
	.zero(gpio4_7_zero)
    );

    sky130_ef_io__gpiov2_pad gpio8_0_pad (
	.IN_H(gpio8_0_in_h),
	.IN(gpio8_0_in),
	.OUT(gpio8_0_out),
	.OE_N(gpio8_0_oe_n),
	.HLD_H_N(gpio8_0_hld_h_n),
	.ENABLE_H(gpio8_0_enable_h),
	.ENABLE_INP_H(gpio8_0_enable_inp_h),
	.ENABLE_VDDA_H(gpio8_0_enable_vdda_h),
	.ENABLE_VDDIO(gpio8_0_enable_vddio),
	.ENABLE_VSWITCH_H(gpio8_0_enable_vswitch_h),
	.INP_DIS(gpio8_0_inp_dis),
	.VTRIP_SEL(gpio8_0_vtrip_sel),
	.SLOW(gpio8_0_slow),
	.HLD_OVR(gpio8_0_hld_ovr),
	.ANALOG_EN(gpio8_0_analog_en),
	.ANALOG_SEL(gpio8_0_analog_sel),
	.ANALOG_POL(gpio8_0_analog_pol),
	.DM(gpio8_0_dm),
	.IB_MODE_SEL(gpio8_0_ib_mode_sel),
	.PAD(gpio8_0),
	.PAD_A_NOESD_H(gpio8_0_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio8_0_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio8_0_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio8_0_tie_hi_esd),
	.TIE_LO_ESD(gpio8_0_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio8_0_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio8_0_one),
	.zero(gpio8_0_zero)
    );

    sky130_ef_io__vdda_hvc_clamped_pad vdda0_0_pad (
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VDDA_PAD(vdda0_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_fd_io__top_gpio_ovtv2 gpio1_4_pad (
	.OUT(gpio1_4_out),
	.OE_N(gpio1_4_oe_n),
	.HLD_H_N(gpio1_4_hld_h_n),
	.ENABLE_H(gpio1_4_enable_h),
	.ENABLE_INP_H(gpio1_4_enable_inp_h),
	.ENABLE_VDDA_H(gpio1_4_enable_vdda_h),
	.ENABLE_VDDIO(gpio1_4_enable_vddio),
	.ENABLE_VSWITCH_H(gpio1_4_enable_vswitch_h),
	.INP_DIS(gpio1_4_inp_dis),
	.VTRIP_SEL(gpio1_4_vtrip_sel),
	.HYS_TRIM(gpio1_4_hys_trim),
	.SLOW(gpio1_4_slow),
	.SLEW_CTL(gpio1_4_slew_ctl),
	.HLD_OVR(gpio1_4_hld_ovr),
	.ANALOG_EN(gpio1_4_analog_en),
	.ANALOG_SEL(gpio1_4_analog_sel),
	.ANALOG_POL(gpio1_4_analog_pol),
	.DM(gpio1_4_dm),
	.IB_MODE_SEL(gpio1_4_ib_mode_sel),
	.VINREF(vref_e_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda1),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio1_4),
	.PAD_A_NOESD_H(gpio1_4_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio1_4_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio1_4_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.IN(gpio1_4_in),
	.IN_H(gpio1_4_in_h),
	.TIE_HI_ESD(gpio1_4_tie_hi_esd),
	.TIE_LO_ESD(gpio1_4_tie_lo_esd)
    );

    constant_block gpio1_4_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio1_4_one),
	.zero(gpio1_4_zero)
    );

    sky130_ef_io__vssio_hvc_clamped_pad vssio_6_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VSSIO_PAD(vssio_6),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio3_7_pad (
	.IN_H(gpio3_7_in_h),
	.IN(gpio3_7_in),
	.OUT(gpio3_7_out),
	.OE_N(gpio3_7_oe_n),
	.HLD_H_N(gpio3_7_hld_h_n),
	.ENABLE_H(gpio3_7_enable_h),
	.ENABLE_INP_H(gpio3_7_enable_inp_h),
	.ENABLE_VDDA_H(gpio3_7_enable_vdda_h),
	.ENABLE_VDDIO(gpio3_7_enable_vddio),
	.ENABLE_VSWITCH_H(gpio3_7_enable_vswitch_h),
	.INP_DIS(gpio3_7_inp_dis),
	.VTRIP_SEL(gpio3_7_vtrip_sel),
	.SLOW(gpio3_7_slow),
	.HLD_OVR(gpio3_7_hld_ovr),
	.ANALOG_EN(gpio3_7_analog_en),
	.ANALOG_SEL(gpio3_7_analog_sel),
	.ANALOG_POL(gpio3_7_analog_pol),
	.DM(gpio3_7_dm),
	.IB_MODE_SEL(gpio3_7_ib_mode_sel),
	.PAD(gpio3_7),
	.PAD_A_NOESD_H(gpio3_7_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio3_7_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio3_7_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio3_7_tie_hi_esd),
	.TIE_LO_ESD(gpio3_7_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio3_7_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio3_7_one),
	.zero(gpio3_7_zero)
    );

    sky130_ef_io__vccd_lvc_clamped3_pad vccd2_0_pad (
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD_PAD(vccd2_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio),
	.VCCD1(vccd2[1]),
	.VSSD1(vssd2[1])
    );

    sky130_ef_io__gpiov2_pad gpio7_0_pad (
	.IN_H(gpio7_0_in_h),
	.IN(gpio7_0_in),
	.OUT(gpio7_0_out),
	.OE_N(gpio7_0_oe_n),
	.HLD_H_N(gpio7_0_hld_h_n),
	.ENABLE_H(gpio7_0_enable_h),
	.ENABLE_INP_H(gpio7_0_enable_inp_h),
	.ENABLE_VDDA_H(gpio7_0_enable_vdda_h),
	.ENABLE_VDDIO(gpio7_0_enable_vddio),
	.ENABLE_VSWITCH_H(gpio7_0_enable_vswitch_h),
	.INP_DIS(gpio7_0_inp_dis),
	.VTRIP_SEL(gpio7_0_vtrip_sel),
	.SLOW(gpio7_0_slow),
	.HLD_OVR(gpio7_0_hld_ovr),
	.ANALOG_EN(gpio7_0_analog_en),
	.ANALOG_SEL(gpio7_0_analog_sel),
	.ANALOG_POL(gpio7_0_analog_pol),
	.DM(gpio7_0_dm),
	.IB_MODE_SEL(gpio7_0_ib_mode_sel),
	.PAD(gpio7_0),
	.PAD_A_NOESD_H(gpio7_0_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio7_0_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio7_0_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio7_0_tie_hi_esd),
	.TIE_LO_ESD(gpio7_0_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio7_0_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio7_0_one),
	.zero(gpio7_0_zero)
    );

    sky130_ef_io__vddio_hvc_clamped_pad vddio_7_pad (
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VDDIO_PAD(vddio_7),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio0_4_pad (
	.IN_H(gpio0_4_in_h),
	.IN(gpio0_4_in),
	.OUT(gpio0_4_out),
	.OE_N(gpio0_4_oe_n),
	.HLD_H_N(gpio0_4_hld_h_n),
	.ENABLE_H(gpio0_4_enable_h),
	.ENABLE_INP_H(gpio0_4_enable_inp_h),
	.ENABLE_VDDA_H(gpio0_4_enable_vdda_h),
	.ENABLE_VDDIO(gpio0_4_enable_vddio),
	.ENABLE_VSWITCH_H(gpio0_4_enable_vswitch_h),
	.INP_DIS(gpio0_4_inp_dis),
	.VTRIP_SEL(gpio0_4_vtrip_sel),
	.SLOW(gpio0_4_slow),
	.HLD_OVR(gpio0_4_hld_ovr),
	.ANALOG_EN(gpio0_4_analog_en),
	.ANALOG_SEL(gpio0_4_analog_sel),
	.ANALOG_POL(gpio0_4_analog_pol),
	.DM(gpio0_4_dm),
	.IB_MODE_SEL(gpio0_4_ib_mode_sel),
	.PAD(gpio0_4),
	.PAD_A_NOESD_H(gpio0_4_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio0_4_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio0_4_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio0_4_tie_hi_esd),
	.TIE_LO_ESD(gpio0_4_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio0_4_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio0_4_one),
	.zero(gpio0_4_zero)
    );

    sky130_ef_io__gpiov2_pad gpio2_7_pad (
	.IN_H(gpio2_7_in_h),
	.IN(gpio2_7_in),
	.OUT(gpio2_7_out),
	.OE_N(gpio2_7_oe_n),
	.HLD_H_N(gpio2_7_hld_h_n),
	.ENABLE_H(gpio2_7_enable_h),
	.ENABLE_INP_H(gpio2_7_enable_inp_h),
	.ENABLE_VDDA_H(gpio2_7_enable_vdda_h),
	.ENABLE_VDDIO(gpio2_7_enable_vddio),
	.ENABLE_VSWITCH_H(gpio2_7_enable_vswitch_h),
	.INP_DIS(gpio2_7_inp_dis),
	.VTRIP_SEL(gpio2_7_vtrip_sel),
	.SLOW(gpio2_7_slow),
	.HLD_OVR(gpio2_7_hld_ovr),
	.ANALOG_EN(gpio2_7_analog_en),
	.ANALOG_SEL(gpio2_7_analog_sel),
	.ANALOG_POL(gpio2_7_analog_pol),
	.DM(gpio2_7_dm),
	.IB_MODE_SEL(gpio2_7_ib_mode_sel),
	.PAD(gpio2_7),
	.PAD_A_NOESD_H(gpio2_7_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio2_7_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio2_7_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio2_7_tie_hi_esd),
	.TIE_LO_ESD(gpio2_7_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio2_7_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio2_7_one),
	.zero(gpio2_7_zero)
    );

    sky130_ef_io__vccd_lvc_clamped3_pad vccd1_0_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD_PAD(vccd1_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio),
	.VCCD1(vccd1[1]),
	.VSSD1(vssd1[1])
    );

    sky130_fd_io__top_gpio_ovtv2 gpio6_0_pad (
	.OUT(gpio6_0_out),
	.OE_N(gpio6_0_oe_n),
	.HLD_H_N(gpio6_0_hld_h_n),
	.ENABLE_H(gpio6_0_enable_h),
	.ENABLE_INP_H(gpio6_0_enable_inp_h),
	.ENABLE_VDDA_H(gpio6_0_enable_vdda_h),
	.ENABLE_VDDIO(gpio6_0_enable_vddio),
	.ENABLE_VSWITCH_H(gpio6_0_enable_vswitch_h),
	.INP_DIS(gpio6_0_inp_dis),
	.VTRIP_SEL(gpio6_0_vtrip_sel),
	.HYS_TRIM(gpio6_0_hys_trim),
	.SLOW(gpio6_0_slow),
	.SLEW_CTL(gpio6_0_slew_ctl),
	.HLD_OVR(gpio6_0_hld_ovr),
	.ANALOG_EN(gpio6_0_analog_en),
	.ANALOG_SEL(gpio6_0_analog_sel),
	.ANALOG_POL(gpio6_0_analog_pol),
	.DM(gpio6_0_dm),
	.IB_MODE_SEL(gpio6_0_ib_mode_sel),
	.VINREF(vref_w_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda2),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio6_0),
	.PAD_A_NOESD_H(gpio6_0_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio6_0_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio6_0_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.IN(gpio6_0_in),
	.IN_H(gpio6_0_in_h),
	.TIE_HI_ESD(gpio6_0_tie_hi_esd),
	.TIE_LO_ESD(gpio6_0_tie_lo_esd)
    );

    constant_block gpio6_0_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio6_0_one),
	.zero(gpio6_0_zero)
    );

    sky130_ef_io__gpiov2_pad gpio8_3_pad (
	.IN_H(gpio8_3_in_h),
	.IN(gpio8_3_in),
	.OUT(gpio8_3_out),
	.OE_N(gpio8_3_oe_n),
	.HLD_H_N(gpio8_3_hld_h_n),
	.ENABLE_H(gpio8_3_enable_h),
	.ENABLE_INP_H(gpio8_3_enable_inp_h),
	.ENABLE_VDDA_H(gpio8_3_enable_vdda_h),
	.ENABLE_VDDIO(gpio8_3_enable_vddio),
	.ENABLE_VSWITCH_H(gpio8_3_enable_vswitch_h),
	.INP_DIS(gpio8_3_inp_dis),
	.VTRIP_SEL(gpio8_3_vtrip_sel),
	.SLOW(gpio8_3_slow),
	.HLD_OVR(gpio8_3_hld_ovr),
	.ANALOG_EN(gpio8_3_analog_en),
	.ANALOG_SEL(gpio8_3_analog_sel),
	.ANALOG_POL(gpio8_3_analog_pol),
	.DM(gpio8_3_dm),
	.IB_MODE_SEL(gpio8_3_ib_mode_sel),
	.PAD(gpio8_3),
	.PAD_A_NOESD_H(gpio8_3_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio8_3_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio8_3_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio8_3_tie_hi_esd),
	.TIE_LO_ESD(gpio8_3_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio8_3_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio8_3_one),
	.zero(gpio8_3_zero)
    );

    sky130_fd_io__top_analog_pad xo1_pad (
	.pad_core(xo1_core),
	.pad(xo1),
	.amuxbus_a(amuxbus_a_s),
	.amuxbus_b(amuxbus_b_s),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda3),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa3),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio)
    );

    sky130_fd_io__top_gpio_ovtv2 gpio1_7_pad (
	.OUT(gpio1_7_out),
	.OE_N(gpio1_7_oe_n),
	.HLD_H_N(gpio1_7_hld_h_n),
	.ENABLE_H(gpio1_7_enable_h),
	.ENABLE_INP_H(gpio1_7_enable_inp_h),
	.ENABLE_VDDA_H(gpio1_7_enable_vdda_h),
	.ENABLE_VDDIO(gpio1_7_enable_vddio),
	.ENABLE_VSWITCH_H(gpio1_7_enable_vswitch_h),
	.INP_DIS(gpio1_7_inp_dis),
	.VTRIP_SEL(gpio1_7_vtrip_sel),
	.HYS_TRIM(gpio1_7_hys_trim),
	.SLOW(gpio1_7_slow),
	.SLEW_CTL(gpio1_7_slew_ctl),
	.HLD_OVR(gpio1_7_hld_ovr),
	.ANALOG_EN(gpio1_7_analog_en),
	.ANALOG_SEL(gpio1_7_analog_sel),
	.ANALOG_POL(gpio1_7_analog_pol),
	.DM(gpio1_7_dm),
	.IB_MODE_SEL(gpio1_7_ib_mode_sel),
	.VINREF(vref_e_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda1),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio1_7),
	.PAD_A_NOESD_H(gpio1_7_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio1_7_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio1_7_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.IN(gpio1_7_in),
	.IN_H(gpio1_7_in_h),
	.TIE_HI_ESD(gpio1_7_tie_hi_esd),
	.TIE_LO_ESD(gpio1_7_tie_lo_esd)
    );

    constant_block gpio1_7_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio1_7_one),
	.zero(gpio1_7_zero)
    );

    sky130_ef_io__vccd_lvc_clamped_pad vccd0_0_pad (
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VCCD_PAD(vccd0_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio5_0_pad (
	.IN_H(gpio5_0_in_h),
	.IN(gpio5_0_in),
	.OUT(gpio5_0_out),
	.OE_N(gpio5_0_oe_n),
	.HLD_H_N(gpio5_0_hld_h_n),
	.ENABLE_H(gpio5_0_enable_h),
	.ENABLE_INP_H(gpio5_0_enable_inp_h),
	.ENABLE_VDDA_H(gpio5_0_enable_vdda_h),
	.ENABLE_VDDIO(gpio5_0_enable_vddio),
	.ENABLE_VSWITCH_H(gpio5_0_enable_vswitch_h),
	.INP_DIS(gpio5_0_inp_dis),
	.VTRIP_SEL(gpio5_0_vtrip_sel),
	.SLOW(gpio5_0_slow),
	.HLD_OVR(gpio5_0_hld_ovr),
	.ANALOG_EN(gpio5_0_analog_en),
	.ANALOG_SEL(gpio5_0_analog_sel),
	.ANALOG_POL(gpio5_0_analog_pol),
	.DM(gpio5_0_dm),
	.IB_MODE_SEL(gpio5_0_ib_mode_sel),
	.PAD(gpio5_0),
	.PAD_A_NOESD_H(gpio5_0_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio5_0_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio5_0_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio5_0_tie_hi_esd),
	.TIE_LO_ESD(gpio5_0_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio5_0_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio5_0_one),
	.zero(gpio5_0_zero)
    );

    sky130_fd_io__top_vrefcapv2 vcap_w (
	.amuxbus_a(amuxbus_a_w),
	.amuxbus_b(amuxbus_b_w),
	.cneg(vssio_q),
	.cpos(vref_w_vinref),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda2),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa2),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio)
    );

    sky130_ef_io__vssio_hvc_clamped_pad vssio_9_pad (
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VSSIO_PAD(vssio_9),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio7_3_pad (
	.IN_H(gpio7_3_in_h),
	.IN(gpio7_3_in),
	.OUT(gpio7_3_out),
	.OE_N(gpio7_3_oe_n),
	.HLD_H_N(gpio7_3_hld_h_n),
	.ENABLE_H(gpio7_3_enable_h),
	.ENABLE_INP_H(gpio7_3_enable_inp_h),
	.ENABLE_VDDA_H(gpio7_3_enable_vdda_h),
	.ENABLE_VDDIO(gpio7_3_enable_vddio),
	.ENABLE_VSWITCH_H(gpio7_3_enable_vswitch_h),
	.INP_DIS(gpio7_3_inp_dis),
	.VTRIP_SEL(gpio7_3_vtrip_sel),
	.SLOW(gpio7_3_slow),
	.HLD_OVR(gpio7_3_hld_ovr),
	.ANALOG_EN(gpio7_3_analog_en),
	.ANALOG_SEL(gpio7_3_analog_sel),
	.ANALOG_POL(gpio7_3_analog_pol),
	.DM(gpio7_3_dm),
	.IB_MODE_SEL(gpio7_3_ib_mode_sel),
	.PAD(gpio7_3),
	.PAD_A_NOESD_H(gpio7_3_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio7_3_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio7_3_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio7_3_tie_hi_esd),
	.TIE_LO_ESD(gpio7_3_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio7_3_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio7_3_one),
	.zero(gpio7_3_zero)
    );

    sky130_ef_io__gpiov2_pad gpio0_7_pad (
	.IN_H(gpio0_7_in_h),
	.IN(gpio0_7_in),
	.OUT(gpio0_7_out),
	.OE_N(gpio0_7_oe_n),
	.HLD_H_N(gpio0_7_hld_h_n),
	.ENABLE_H(gpio0_7_enable_h),
	.ENABLE_INP_H(gpio0_7_enable_inp_h),
	.ENABLE_VDDA_H(gpio0_7_enable_vdda_h),
	.ENABLE_VDDIO(gpio0_7_enable_vddio),
	.ENABLE_VSWITCH_H(gpio0_7_enable_vswitch_h),
	.INP_DIS(gpio0_7_inp_dis),
	.VTRIP_SEL(gpio0_7_vtrip_sel),
	.SLOW(gpio0_7_slow),
	.HLD_OVR(gpio0_7_hld_ovr),
	.ANALOG_EN(gpio0_7_analog_en),
	.ANALOG_SEL(gpio0_7_analog_sel),
	.ANALOG_POL(gpio0_7_analog_pol),
	.DM(gpio0_7_dm),
	.IB_MODE_SEL(gpio0_7_ib_mode_sel),
	.PAD(gpio0_7),
	.PAD_A_NOESD_H(gpio0_7_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio0_7_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio0_7_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio0_7_tie_hi_esd),
	.TIE_LO_ESD(gpio0_7_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio0_7_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio0_7_one),
	.zero(gpio0_7_zero)
    );

    sky130_ef_io__gpiov2_pad gpio4_0_pad (
	.IN_H(gpio4_0_in_h),
	.IN(gpio4_0_in),
	.OUT(gpio4_0_out),
	.OE_N(gpio4_0_oe_n),
	.HLD_H_N(gpio4_0_hld_h_n),
	.ENABLE_H(gpio4_0_enable_h),
	.ENABLE_INP_H(gpio4_0_enable_inp_h),
	.ENABLE_VDDA_H(gpio4_0_enable_vdda_h),
	.ENABLE_VDDIO(gpio4_0_enable_vddio),
	.ENABLE_VSWITCH_H(gpio4_0_enable_vswitch_h),
	.INP_DIS(gpio4_0_inp_dis),
	.VTRIP_SEL(gpio4_0_vtrip_sel),
	.SLOW(gpio4_0_slow),
	.HLD_OVR(gpio4_0_hld_ovr),
	.ANALOG_EN(gpio4_0_analog_en),
	.ANALOG_SEL(gpio4_0_analog_sel),
	.ANALOG_POL(gpio4_0_analog_pol),
	.DM(gpio4_0_dm),
	.IB_MODE_SEL(gpio4_0_ib_mode_sel),
	.PAD(gpio4_0),
	.PAD_A_NOESD_H(gpio4_0_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio4_0_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio4_0_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio4_0_tie_hi_esd),
	.TIE_LO_ESD(gpio4_0_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio4_0_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio4_0_one),
	.zero(gpio4_0_zero)
    );

    sky130_fd_io__top_gpio_ovtv2 gpio6_3_pad (
	.OUT(gpio6_3_out),
	.OE_N(gpio6_3_oe_n),
	.HLD_H_N(gpio6_3_hld_h_n),
	.ENABLE_H(gpio6_3_enable_h),
	.ENABLE_INP_H(gpio6_3_enable_inp_h),
	.ENABLE_VDDA_H(gpio6_3_enable_vdda_h),
	.ENABLE_VDDIO(gpio6_3_enable_vddio),
	.ENABLE_VSWITCH_H(gpio6_3_enable_vswitch_h),
	.INP_DIS(gpio6_3_inp_dis),
	.VTRIP_SEL(gpio6_3_vtrip_sel),
	.HYS_TRIM(gpio6_3_hys_trim),
	.SLOW(gpio6_3_slow),
	.SLEW_CTL(gpio6_3_slew_ctl),
	.HLD_OVR(gpio6_3_hld_ovr),
	.ANALOG_EN(gpio6_3_analog_en),
	.ANALOG_SEL(gpio6_3_analog_sel),
	.ANALOG_POL(gpio6_3_analog_pol),
	.DM(gpio6_3_dm),
	.IB_MODE_SEL(gpio6_3_ib_mode_sel),
	.VINREF(vref_w_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda2),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio6_3),
	.PAD_A_NOESD_H(gpio6_3_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio6_3_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio6_3_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.IN(gpio6_3_in),
	.IN_H(gpio6_3_in_h),
	.TIE_HI_ESD(gpio6_3_tie_hi_esd),
	.TIE_LO_ESD(gpio6_3_tie_lo_esd)
    );

    constant_block gpio6_3_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio6_3_one),
	.zero(gpio6_3_zero)
    );

    sky130_ef_io__vssd_lvc_clamped3_pad vssd2_0_pad (
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VSSD_PAD(vssd2_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio),
	.VCCD1(vccd2[0]),
	.VSSD1(vssd2[0])
    );

    sky130_ef_io__gpiov2_pad gpio8_6_pad (
	.IN_H(gpio8_6_in_h),
	.IN(gpio8_6_in),
	.OUT(gpio8_6_out),
	.OE_N(gpio8_6_oe_n),
	.HLD_H_N(gpio8_6_hld_h_n),
	.ENABLE_H(gpio8_6_enable_h),
	.ENABLE_INP_H(gpio8_6_enable_inp_h),
	.ENABLE_VDDA_H(gpio8_6_enable_vdda_h),
	.ENABLE_VDDIO(gpio8_6_enable_vddio),
	.ENABLE_VSWITCH_H(gpio8_6_enable_vswitch_h),
	.INP_DIS(gpio8_6_inp_dis),
	.VTRIP_SEL(gpio8_6_vtrip_sel),
	.SLOW(gpio8_6_slow),
	.HLD_OVR(gpio8_6_hld_ovr),
	.ANALOG_EN(gpio8_6_analog_en),
	.ANALOG_SEL(gpio8_6_analog_sel),
	.ANALOG_POL(gpio8_6_analog_pol),
	.DM(gpio8_6_dm),
	.IB_MODE_SEL(gpio8_6_ib_mode_sel),
	.PAD(gpio8_6),
	.PAD_A_NOESD_H(gpio8_6_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio8_6_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio8_6_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio8_6_tie_hi_esd),
	.TIE_LO_ESD(gpio8_6_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio8_6_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio8_6_one),
	.zero(gpio8_6_zero)
    );

    sky130_ef_io__gpiov2_pad gpio3_0_pad (
	.IN_H(gpio3_0_in_h),
	.IN(gpio3_0_in),
	.OUT(gpio3_0_out),
	.OE_N(gpio3_0_oe_n),
	.HLD_H_N(gpio3_0_hld_h_n),
	.ENABLE_H(gpio3_0_enable_h),
	.ENABLE_INP_H(gpio3_0_enable_inp_h),
	.ENABLE_VDDA_H(gpio3_0_enable_vdda_h),
	.ENABLE_VDDIO(gpio3_0_enable_vddio),
	.ENABLE_VSWITCH_H(gpio3_0_enable_vswitch_h),
	.INP_DIS(gpio3_0_inp_dis),
	.VTRIP_SEL(gpio3_0_vtrip_sel),
	.SLOW(gpio3_0_slow),
	.HLD_OVR(gpio3_0_hld_ovr),
	.ANALOG_EN(gpio3_0_analog_en),
	.ANALOG_SEL(gpio3_0_analog_sel),
	.ANALOG_POL(gpio3_0_analog_pol),
	.DM(gpio3_0_dm),
	.IB_MODE_SEL(gpio3_0_ib_mode_sel),
	.PAD(gpio3_0),
	.PAD_A_NOESD_H(gpio3_0_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio3_0_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio3_0_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio3_0_tie_hi_esd),
	.TIE_LO_ESD(gpio3_0_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio3_0_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio3_0_one),
	.zero(gpio3_0_zero)
    );

    sky130_ef_io__gpiov2_pad gpio5_3_pad (
	.IN_H(gpio5_3_in_h),
	.IN(gpio5_3_in),
	.OUT(gpio5_3_out),
	.OE_N(gpio5_3_oe_n),
	.HLD_H_N(gpio5_3_hld_h_n),
	.ENABLE_H(gpio5_3_enable_h),
	.ENABLE_INP_H(gpio5_3_enable_inp_h),
	.ENABLE_VDDA_H(gpio5_3_enable_vdda_h),
	.ENABLE_VDDIO(gpio5_3_enable_vddio),
	.ENABLE_VSWITCH_H(gpio5_3_enable_vswitch_h),
	.INP_DIS(gpio5_3_inp_dis),
	.VTRIP_SEL(gpio5_3_vtrip_sel),
	.SLOW(gpio5_3_slow),
	.HLD_OVR(gpio5_3_hld_ovr),
	.ANALOG_EN(gpio5_3_analog_en),
	.ANALOG_SEL(gpio5_3_analog_sel),
	.ANALOG_POL(gpio5_3_analog_pol),
	.DM(gpio5_3_dm),
	.IB_MODE_SEL(gpio5_3_ib_mode_sel),
	.PAD(gpio5_3),
	.PAD_A_NOESD_H(gpio5_3_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio5_3_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio5_3_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio5_3_tie_hi_esd),
	.TIE_LO_ESD(gpio5_3_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio5_3_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio5_3_one),
	.zero(gpio5_3_zero)
    );

    sky130_ef_io__vssd_lvc_clamped3_pad vssd1_0_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VSSD_PAD(vssd1_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio),
	.VCCD1(vccd1[0]),
	.VSSD1(vssd1[0])
    );

    sky130_ef_io__gpiov2_pad gpio7_6_pad (
	.IN_H(gpio7_6_in_h),
	.IN(gpio7_6_in),
	.OUT(gpio7_6_out),
	.OE_N(gpio7_6_oe_n),
	.HLD_H_N(gpio7_6_hld_h_n),
	.ENABLE_H(gpio7_6_enable_h),
	.ENABLE_INP_H(gpio7_6_enable_inp_h),
	.ENABLE_VDDA_H(gpio7_6_enable_vdda_h),
	.ENABLE_VDDIO(gpio7_6_enable_vddio),
	.ENABLE_VSWITCH_H(gpio7_6_enable_vswitch_h),
	.INP_DIS(gpio7_6_inp_dis),
	.VTRIP_SEL(gpio7_6_vtrip_sel),
	.SLOW(gpio7_6_slow),
	.HLD_OVR(gpio7_6_hld_ovr),
	.ANALOG_EN(gpio7_6_analog_en),
	.ANALOG_SEL(gpio7_6_analog_sel),
	.ANALOG_POL(gpio7_6_analog_pol),
	.DM(gpio7_6_dm),
	.IB_MODE_SEL(gpio7_6_ib_mode_sel),
	.PAD(gpio7_6),
	.PAD_A_NOESD_H(gpio7_6_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio7_6_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio7_6_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio7_6_tie_hi_esd),
	.TIE_LO_ESD(gpio7_6_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda2),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio7_6_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio7_6_one),
	.zero(gpio7_6_zero)
    );

    sky130_ef_io__vddio_hvc_clamped_pad vddio_0_pad (
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VDDIO_PAD(vddio_0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio2_0_pad (
	.IN_H(gpio2_0_in_h),
	.IN(gpio2_0_in),
	.OUT(gpio2_0_out),
	.OE_N(gpio2_0_oe_n),
	.HLD_H_N(gpio2_0_hld_h_n),
	.ENABLE_H(gpio2_0_enable_h),
	.ENABLE_INP_H(gpio2_0_enable_inp_h),
	.ENABLE_VDDA_H(gpio2_0_enable_vdda_h),
	.ENABLE_VDDIO(gpio2_0_enable_vddio),
	.ENABLE_VSWITCH_H(gpio2_0_enable_vswitch_h),
	.INP_DIS(gpio2_0_inp_dis),
	.VTRIP_SEL(gpio2_0_vtrip_sel),
	.SLOW(gpio2_0_slow),
	.HLD_OVR(gpio2_0_hld_ovr),
	.ANALOG_EN(gpio2_0_analog_en),
	.ANALOG_SEL(gpio2_0_analog_sel),
	.ANALOG_POL(gpio2_0_analog_pol),
	.DM(gpio2_0_dm),
	.IB_MODE_SEL(gpio2_0_ib_mode_sel),
	.PAD(gpio2_0),
	.PAD_A_NOESD_H(gpio2_0_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio2_0_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio2_0_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio2_0_tie_hi_esd),
	.TIE_LO_ESD(gpio2_0_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_e),
	.AMUXBUS_B(amuxbus_b_e),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda1),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa1),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio2_0_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio2_0_one),
	.zero(gpio2_0_zero)
    );

    sky130_fd_io__top_analog_pad analog_1_pad (
	.pad_core(analog_1_core),
	.pad(analog_1),
	.amuxbus_a(amuxbus_a_n),
	.amuxbus_b(amuxbus_b_n),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda0),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa0),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio)
    );

    sky130_ef_io__vssd_lvc_clamped_pad vssd0_0_pad (
	.AMUXBUS_A(amuxbus_a_s),
	.AMUXBUS_B(amuxbus_b_s),
	.VSSD_PAD(vssd0_0),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda3),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa3),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    sky130_ef_io__gpiov2_pad gpio4_3_pad (
	.IN_H(gpio4_3_in_h),
	.IN(gpio4_3_in),
	.OUT(gpio4_3_out),
	.OE_N(gpio4_3_oe_n),
	.HLD_H_N(gpio4_3_hld_h_n),
	.ENABLE_H(gpio4_3_enable_h),
	.ENABLE_INP_H(gpio4_3_enable_inp_h),
	.ENABLE_VDDA_H(gpio4_3_enable_vdda_h),
	.ENABLE_VDDIO(gpio4_3_enable_vddio),
	.ENABLE_VSWITCH_H(gpio4_3_enable_vswitch_h),
	.INP_DIS(gpio4_3_inp_dis),
	.VTRIP_SEL(gpio4_3_vtrip_sel),
	.SLOW(gpio4_3_slow),
	.HLD_OVR(gpio4_3_hld_ovr),
	.ANALOG_EN(gpio4_3_analog_en),
	.ANALOG_SEL(gpio4_3_analog_sel),
	.ANALOG_POL(gpio4_3_analog_pol),
	.DM(gpio4_3_dm),
	.IB_MODE_SEL(gpio4_3_ib_mode_sel),
	.PAD(gpio4_3),
	.PAD_A_NOESD_H(gpio4_3_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio4_3_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio4_3_pad_a_esd_1_h),
	.TIE_HI_ESD(gpio4_3_tie_hi_esd),
	.TIE_LO_ESD(gpio4_3_tie_lo_esd),
	.AMUXBUS_A(amuxbus_a_n),
	.AMUXBUS_B(amuxbus_b_n),
	.VCCD(vccd0),
	.VCCHIB(vccd0),
	.VDDA(vdda0),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VSSA(vssa0),
	.VSSD(vssd0),
	.VSSIO(vssio),
	.VSSIO_Q(vssio_q),
	.VSWITCH(vddio)
    );

    constant_block gpio4_3_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio4_3_one),
	.zero(gpio4_3_zero)
    );

    sky130_fd_io__top_gpio_ovtv2 gpio6_6_pad (
	.OUT(gpio6_6_out),
	.OE_N(gpio6_6_oe_n),
	.HLD_H_N(gpio6_6_hld_h_n),
	.ENABLE_H(gpio6_6_enable_h),
	.ENABLE_INP_H(gpio6_6_enable_inp_h),
	.ENABLE_VDDA_H(gpio6_6_enable_vdda_h),
	.ENABLE_VDDIO(gpio6_6_enable_vddio),
	.ENABLE_VSWITCH_H(gpio6_6_enable_vswitch_h),
	.INP_DIS(gpio6_6_inp_dis),
	.VTRIP_SEL(gpio6_6_vtrip_sel),
	.HYS_TRIM(gpio6_6_hys_trim),
	.SLOW(gpio6_6_slow),
	.SLEW_CTL(gpio6_6_slew_ctl),
	.HLD_OVR(gpio6_6_hld_ovr),
	.ANALOG_EN(gpio6_6_analog_en),
	.ANALOG_SEL(gpio6_6_analog_sel),
	.ANALOG_POL(gpio6_6_analog_pol),
	.DM(gpio6_6_dm),
	.IB_MODE_SEL(gpio6_6_ib_mode_sel),
	.VINREF(vref_w_vinref),
	.VDDIO(vddio),
	.VDDIO_Q(vddio_q),
	.VDDA(vdda2),
	.VCCD(vccd0),
	.VSWITCH(vddio),
	.VCCHIB(vccd0),
	.VSSA(vssa2),
	.VSSD(vssd0),
	.VSSIO_Q(vssio_q),
	.VSSIO(vssio),
	.PAD(gpio6_6),
	.PAD_A_NOESD_H(gpio6_6_pad_a_noesd_h),
	.PAD_A_ESD_0_H(gpio6_6_pad_a_esd_0_h),
	.PAD_A_ESD_1_H(gpio6_6_pad_a_esd_1_h),
	.AMUXBUS_A(amuxbus_a_w),
	.AMUXBUS_B(amuxbus_b_w),
	.IN(gpio6_6_in),
	.IN_H(gpio6_6_in_h),
	.TIE_HI_ESD(gpio6_6_tie_hi_esd),
	.TIE_LO_ESD(gpio6_6_tie_lo_esd)
    );

    constant_block gpio6_6_const (
	.vccd(vccd0),
	.vssd(vssd0),
	.one(gpio6_6_one),
	.zero(gpio6_6_zero)
    );

    sky130_fd_io__top_analog_pad xi0_pad (
	.pad_core(xi0_core),
	.pad(xi0),
	.amuxbus_a(amuxbus_a_s),
	.amuxbus_b(amuxbus_b_s),
	.vccd(vccd0),
	.vcchib(vccd0),
	.vdda(vdda3),
	.vddio(vddio),
	.vddio_q(vddio_q),
	.vssa(vssa3),
	.vssd(vssd0),
	.vssio(vssio),
	.vssio_q(vssio_q),
	.vswitch(vddio)
    );

    /* Additional modules */
    /* Level shifted output for the RESETB pin */

    xres_lvlshift xres_lvlshift_0 (
    `ifdef USE_POWER_PINS
	.VPWR(vddio),
	.VGND(vssio),
	.LVPWR(vccd0),
	.LVGND(vssd0),
    `endif
	.A(resetb_xres_h_n),
	.X(resetb_xres_n)
    );

    /* Product ID (note:  Unprogrammed version) */
    product_id_rom_8bit product_id_rom_8bit_0 (
    `ifdef USE_POWER_PINS
	.VPWR(vccd),
	.VGND(vssd),
    `endif
	.product_id(product_id)
    );

    /* Project (user) ID (note:  Unprogrammed version) */
    project_id_rom_32bit project_id_rom_32bit_0 (
    `ifdef USE_POWER_PINS
	.VPWR(vccd),
	.VGND(vssd),
    `endif
	.project_id(project_id)
    );

endmodule

`default_nettype wire
