magic
tech sky130A
magscale 1 2
timestamp 1726510490
<< checkpaint >>
rect -1205 8088 1531 14399
rect -1212 4792 1531 8088
rect -1212 4721 1503 4792
<< metal2 >>
rect 75 13132 85 13134
rect 0 13080 85 13132
rect 75 13078 85 13080
rect 255 13078 264 13134
rect 75 12151 85 12153
rect 0 12099 85 12151
rect 75 12097 85 12099
rect 255 12097 264 12153
rect 0 7620 264 7625
rect 0 7502 85 7620
rect 255 7502 264 7620
rect 0 7497 264 7502
rect 75 6797 85 6799
rect 0 6745 85 6797
rect 75 6743 85 6745
rect 255 6743 264 6799
rect 75 6599 85 6601
rect 0 6547 85 6599
rect 75 6545 85 6547
rect 255 6545 264 6601
rect 75 6399 85 6401
rect 0 6347 85 6399
rect 75 6345 85 6347
rect 255 6345 264 6401
rect 75 6111 85 6113
rect 0 6059 85 6111
rect 75 6057 85 6059
rect 255 6057 264 6113
rect 60 1283 70 1285
rect 0 1231 70 1283
rect 60 1229 70 1231
rect 240 1229 249 1285
rect 60 1031 70 1033
rect 0 979 70 1031
rect 60 977 70 979
rect 240 977 249 1033
<< via2 >>
rect 85 13078 255 13134
rect 85 12097 255 12153
rect 85 7502 255 7620
rect 85 6743 255 6799
rect 85 6545 255 6601
rect 85 6345 255 6401
rect 85 6057 255 6113
rect 70 1229 240 1285
rect 70 977 240 1033
<< metal3 >>
rect 80 13136 260 13139
rect 80 13134 300 13136
rect 80 13078 85 13134
rect 255 13078 300 13134
rect 80 13076 300 13078
rect 80 13073 260 13076
rect 80 12155 260 12158
rect 80 12153 300 12155
rect 80 12097 85 12153
rect 255 12097 300 12153
rect 80 12095 300 12097
rect 80 12092 260 12095
rect 80 7620 300 7625
rect 80 7502 85 7620
rect 255 7502 300 7620
rect 80 7497 300 7502
rect 80 6801 260 6804
rect 80 6799 300 6801
rect 80 6743 85 6799
rect 255 6743 300 6799
rect 80 6741 300 6743
rect 80 6738 260 6741
rect 80 6603 260 6606
rect 80 6601 300 6603
rect 80 6545 85 6601
rect 255 6545 300 6601
rect 80 6543 300 6545
rect 80 6540 260 6543
rect 80 6403 260 6406
rect 80 6401 300 6403
rect 80 6345 85 6401
rect 255 6345 300 6401
rect 80 6343 300 6345
rect 80 6340 260 6343
rect 80 6115 260 6118
rect 80 6113 300 6115
rect 80 6057 85 6113
rect 255 6057 300 6113
rect 80 6055 300 6057
rect 80 6052 260 6055
rect 65 1287 245 1290
rect 65 1285 300 1287
rect 65 1229 70 1285
rect 240 1229 300 1285
rect 65 1227 300 1229
rect 65 1224 245 1227
rect 65 1035 245 1038
rect 65 1033 300 1035
rect 65 977 70 1033
rect 240 977 300 1033
rect 65 975 300 977
rect 65 972 245 975
<< labels >>
flabel metal3 s 240 12095 300 12155 0 FreeSans 480 0 0 0 ref_sel<0>
port 5 nsew
flabel metal3 s 240 13076 300 13136 0 FreeSans 480 0 0 0 ref_sel<1>
port 6 nsew
flabel metal3 s 240 7497 300 7625 0 FreeSans 480 0 0 0 vinref
port 7 nsew
flabel metal3 s 240 975 300 1035 0 FreeSans 480 0 0 0 ref_sel<3>
port 8 nsew
flabel metal3 s 240 1227 300 1287 0 FreeSans 480 0 0 0 ref_sel<4>
port 9 nsew
flabel metal3 s 240 6741 300 6801 0 FreeSans 480 0 0 0 ref_sel<2>
port 4 nsew
flabel metal3 s 240 6543 300 6603 0 FreeSans 480 0 0 0 enable_h
port 3 nsew
flabel metal3 s 240 6343 300 6403 0 FreeSans 480 0 0 0 hld_h_n
port 2 nsew
flabel metal3 s 240 6055 300 6115 0 FreeSans 480 0 0 0 vrefgen_en
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 300 16000
string flatten true
<< end >>
