magic
tech sky130A
magscale 1 2
timestamp 1719074309
<< metal2 >>
rect 60 7210 70 7212
rect 0 7158 70 7210
rect 60 7156 70 7158
rect 240 7156 250 7212
rect 60 6330 70 6332
rect 0 6278 70 6330
rect 60 6276 70 6278
rect 240 6276 250 6332
rect 60 2708 70 2710
rect 0 2656 70 2708
rect 60 2654 70 2656
rect 240 2654 250 2710
rect 60 2456 70 2458
rect 0 2404 70 2456
rect 60 2402 70 2404
rect 240 2402 250 2458
rect 60 2204 70 2206
rect 0 2152 70 2204
rect 60 2150 70 2152
rect 240 2150 250 2206
rect 60 1952 70 1954
rect 0 1900 70 1952
rect 60 1898 70 1900
rect 240 1898 250 1954
rect 60 1700 70 1702
rect 0 1648 70 1700
rect 60 1646 70 1648
rect 240 1646 250 1702
rect 60 1364 70 1366
rect 0 1312 70 1364
rect 60 1310 70 1312
rect 240 1310 250 1366
<< via2 >>
rect 70 7156 240 7212
rect 70 6276 240 6332
rect 70 2654 240 2710
rect 70 2402 240 2458
rect 70 2150 240 2206
rect 70 1898 240 1954
rect 70 1646 240 1702
rect 70 1310 240 1366
<< metal3 >>
rect 65 7214 245 7217
rect 65 7212 300 7214
rect 65 7156 70 7212
rect 240 7156 300 7212
rect 65 7154 300 7156
rect 65 7151 245 7154
rect 65 6334 245 6337
rect 65 6332 300 6334
rect 65 6276 70 6332
rect 240 6276 300 6332
rect 65 6274 300 6276
rect 65 6271 245 6274
rect 65 2712 245 2715
rect 65 2710 300 2712
rect 65 2654 70 2710
rect 240 2654 300 2710
rect 65 2652 300 2654
rect 65 2649 245 2652
rect 65 2460 245 2463
rect 65 2458 300 2460
rect 65 2402 70 2458
rect 240 2402 300 2458
rect 65 2400 300 2402
rect 65 2397 245 2400
rect 65 2208 245 2211
rect 65 2206 300 2208
rect 65 2150 70 2206
rect 240 2150 300 2206
rect 65 2148 300 2150
rect 65 2145 245 2148
rect 65 1956 245 1959
rect 65 1954 300 1956
rect 65 1898 70 1954
rect 240 1898 300 1954
rect 65 1896 300 1898
rect 65 1893 245 1896
rect 65 1704 245 1707
rect 65 1702 300 1704
rect 65 1646 70 1702
rect 240 1646 300 1702
rect 65 1644 300 1646
rect 65 1641 245 1644
rect 65 1368 245 1371
rect 65 1366 300 1368
rect 65 1310 70 1366
rect 240 1310 300 1366
rect 65 1308 300 1310
rect 65 1305 245 1308
<< labels >>
flabel metal3 s 240 6274 300 6334 0 FreeSans 480 0 0 0 enable_vdda_h
port 7 nsew
flabel metal3 s 240 7154 300 7214 0 FreeSans 480 0 0 0 hld_vdda_h_n
port 8 nsew
flabel metal3 s 240 2652 300 2712 0 FreeSans 480 0 0 0 switch_aa_sl
port 6 nsew
flabel metal3 s 240 2400 300 2460 0 FreeSans 480 0 0 0 switch_aa_s0
port 5 nsew
flabel metal3 s 240 2148 300 2208 0 FreeSans 480 0 0 0 switch_bb_s0
port 4 nsew
flabel metal3 s 240 1896 300 1956 0 FreeSans 480 0 0 0 switch_bb_sl
port 3 nsew
flabel metal3 s 240 1644 300 1704 0 FreeSans 480 0 0 0 switch_bb_sr
port 2 nsew
flabel metal3 s 240 1308 300 1368 0 FreeSans 480 0 0 0 switch_aa_sr
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 300 9600
string flatten true
<< end >>
