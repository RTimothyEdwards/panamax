magic
tech sky130A
timestamp 1746202547
<< checkpaint >>
rect 1823 4736 6828 5816
rect -302 -326 19590 4736
rect -302 -1384 6538 -326
rect 16420 -398 19300 -326
<< fillblock >>
rect 0 0 17188 4418
use alpha_0  alphaX_0 hexdigits
timestamp 1598786981
transform 1 0 15215 0 1 326
box 0 0 1620 3780
use alpha_0  alphaX_1
timestamp 1598786981
transform 1 0 13078 0 1 326
box 0 0 1620 3780
use alpha_0  alphaX_2
timestamp 1598786981
transform 1 0 10953 0 1 326
box 0 0 1620 3780
use alpha_0  alphaX_3
timestamp 1598786981
transform 1 0 8828 0 1 326
box 0 0 1620 3780
use alpha_0  alphaX_4
timestamp 1598786981
transform 1 0 6703 0 1 326
box 0 0 1620 3780
use alpha_0  alphaX_5
timestamp 1598786981
transform 1 0 4578 0 1 326
box 0 0 1620 3780
use alpha_0  alphaX_6
timestamp 1598786981
transform 1 0 2453 0 1 326
box 0 0 1620 3780
use alpha_0  alphaX_7
timestamp 1598786981
transform 1 0 328 0 1 326
box 0 0 1620 3780
<< end >>
