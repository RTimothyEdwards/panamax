magic
tech sky130A
magscale 1 2
timestamp 1726600167
<< checkpaint >>
rect -1260 998860 718860 1038860
rect -1261 998060 718860 998860
rect -1261 996747 718861 998060
rect -1261 996340 42060 996747
rect -1261 988260 41560 996340
rect 43540 994570 63247 996747
rect 66397 996340 87918 996747
rect 90397 996340 111918 996747
rect 114397 996340 135918 996747
rect 138397 996340 159918 996747
rect 66516 995430 87918 996340
rect 90516 995430 111918 996340
rect 114516 995430 135918 996340
rect 138516 995430 159918 996340
rect 162540 996340 180060 996747
rect 162540 995547 170060 996340
rect 172540 995547 180060 996340
rect 185540 994570 205247 996747
rect 208397 996340 229918 996747
rect 232397 996340 253918 996747
rect 256397 996340 277918 996747
rect 280397 996340 301918 996747
rect 208516 995430 229918 996340
rect 232516 995430 253918 996340
rect 256516 995430 277918 996340
rect 280516 995430 301918 996340
rect 304540 996340 322060 996747
rect 327460 996740 345140 996747
rect 350460 996740 370998 996747
rect 304540 995547 312060 996340
rect 314540 995547 322060 996340
rect 327540 995940 345060 996740
rect 350540 995940 370998 996740
rect 366340 995340 370998 995940
rect 373540 996340 391060 996747
rect 373540 995547 381060 996340
rect 383540 995547 391060 996340
rect 396540 996340 414060 996747
rect 419397 996340 440918 996747
rect 443397 996340 464918 996747
rect 467397 996340 488918 996747
rect 491397 996340 512918 996747
rect 396540 995547 404060 996340
rect 406540 995547 414060 996340
rect 419516 995430 440918 996340
rect 443516 995430 464918 996340
rect 467516 995430 488918 996340
rect 491516 995430 512918 996340
rect 367236 995133 370166 995340
rect 515540 994570 535247 996747
rect 538540 996340 556060 996747
rect 561397 996340 582918 996747
rect 585397 996340 606918 996747
rect 609397 996340 630918 996747
rect 633397 996340 654918 996747
rect 538540 995547 546060 996340
rect 548540 995547 556060 996340
rect 561516 995430 582918 996340
rect 585516 995430 606918 996340
rect 609516 995430 630918 996340
rect 633516 995430 654918 996340
rect 657540 994570 718861 996747
rect 676040 988323 718861 994570
rect -1261 986740 42053 988260
rect 676340 987460 718861 988323
rect -1260 980740 42053 986740
rect 675547 985940 718861 987460
rect -1260 978260 41260 980740
rect 675547 979940 718860 985940
rect -1260 970740 42053 978260
rect 676340 977460 718860 979940
rect -1260 967447 40853 970740
rect 675547 969940 718860 977460
rect -1260 960338 43030 967447
rect 676747 963460 718860 969940
rect -1260 952650 43528 960338
rect -1260 947740 43030 952650
rect -1260 863696 42102 947740
rect 674570 943753 718860 963460
rect 676747 943603 718860 943753
rect 676340 943504 718860 943603
rect -1260 863597 41260 863696
rect -1260 861260 40853 863597
rect -1260 853740 42053 861260
rect 675498 858740 718860 943504
rect -1260 851260 41260 853740
rect 675547 851940 718860 858740
rect -1260 844460 42053 851260
rect 676340 849460 718860 851940
rect -1260 759696 42102 844460
rect 675547 841940 718860 849460
rect 676747 839603 718860 841940
rect 676340 839504 718860 839603
rect -1260 759597 41260 759696
rect -1260 759447 40853 759597
rect -1260 739740 43030 759447
rect 675498 755460 718860 839504
rect -1260 737260 40853 739740
rect -1260 729740 42053 737260
rect 674570 735753 718860 755460
rect 676747 735460 718860 735753
rect -1260 727260 41260 729740
rect 675547 727940 718860 735460
rect -1260 719740 42053 727260
rect 676340 725460 718860 727940
rect -1260 714260 40853 719740
rect 675547 717940 718860 725460
rect -1260 706740 42053 714260
rect 676747 711460 718860 717940
rect -1260 704260 41260 706740
rect -1260 696740 42053 704260
rect 675547 703940 718860 711460
rect 676340 701460 718860 703940
rect -1260 694260 40853 696740
rect -1260 686740 42053 694260
rect 675547 693940 718860 701460
rect 676747 691460 718860 693940
rect -1260 684260 41260 686740
rect -1260 676740 42053 684260
rect 675547 683940 718860 691460
rect 676340 681460 718860 683940
rect -1260 674471 41860 676740
rect -1411 643660 41860 674471
rect 675547 673940 718860 681460
rect 676747 671572 718860 673940
rect -1260 641471 41860 643660
rect -1411 610660 41860 641471
rect -1260 608471 41860 610660
rect -1411 577660 41860 608471
rect -1260 575471 41860 577660
rect -1411 544660 41860 575471
rect -1260 544628 41860 544660
rect 675740 671540 718860 671572
rect 675740 640729 719011 671540
rect 675740 638540 718860 640729
rect 675740 607729 719011 638540
rect 675740 605540 718860 607729
rect 675740 574729 719011 605540
rect 675740 572540 718860 574729
rect -1260 542260 40853 544628
rect -1260 534740 42053 542260
rect 675740 541729 719011 572540
rect 675740 539460 718860 541729
rect -1260 532260 41260 534740
rect -1260 524740 42053 532260
rect 675547 531940 718860 539460
rect 676340 529460 718860 531940
rect -1260 522116 40853 524740
rect -1260 515799 41260 522116
rect 675547 521940 718860 529460
rect 676747 519316 718860 521940
rect -1260 501112 41560 515799
rect 676340 514888 718860 519316
rect -1260 500140 41260 501112
rect 676040 500201 718860 514888
rect -1260 499847 40853 500140
rect -1260 480140 43030 499847
rect 676340 497340 718860 500201
rect 676747 494860 718860 497340
rect -1260 477871 41860 480140
rect -1411 447060 41860 477871
rect 674570 475153 718860 494860
rect 676747 474972 718860 475153
rect -1260 444871 41860 447060
rect -1411 414060 41860 444871
rect -1260 411871 41860 414060
rect -1411 381060 41860 411871
rect -1260 378871 41860 381060
rect -1411 348060 41860 378871
rect -1260 348028 41860 348060
rect 675740 474940 718860 474972
rect 675740 444129 719011 474940
rect 675740 441940 718860 444129
rect 675740 411129 719011 441940
rect 675740 408940 718860 411129
rect 675740 378129 719011 408940
rect 675740 375940 718860 378129
rect -1260 345660 40853 348028
rect -1260 338140 42053 345660
rect 675740 345129 719011 375940
rect 675740 342860 718860 345129
rect -1260 335660 41260 338140
rect -1260 328140 42053 335660
rect 675547 335340 718860 342860
rect 676340 332860 718860 335340
rect -1260 322660 40853 328140
rect 675547 325340 718860 332860
rect -1260 315140 42053 322660
rect 676747 318860 718860 325340
rect -1260 312660 41260 315140
rect -1260 305140 42053 312660
rect 675547 311340 718860 318860
rect 676340 308860 718860 311340
rect -1260 302660 40853 305140
rect -1260 295140 42053 302660
rect 675547 301340 718860 308860
rect 676747 298860 718860 301340
rect -1260 292660 41260 295140
rect -1260 285860 42053 292660
rect 675547 291340 718860 298860
rect 676340 288860 718860 291340
rect -1260 201096 42102 285860
rect 675547 281340 718860 288860
rect 676747 279003 718860 281340
rect 676340 278904 718860 279003
rect -1260 200997 41260 201096
rect -1260 198660 40853 200997
rect -1260 191140 42053 198660
rect 675498 194140 718860 278904
rect -1260 188660 41260 191140
rect -1260 181140 42053 188660
rect 675547 187340 718860 194140
rect 676340 184860 718860 187340
rect -1260 177847 40853 181140
rect -1260 158140 43030 177847
rect 675547 177340 718860 184860
rect 676747 174860 718860 177340
rect -1260 74096 42102 158140
rect 674570 155153 718860 174860
rect 676747 155003 718860 155153
rect 676340 154904 718860 155003
rect -1260 73997 41260 74096
rect -1260 71660 40853 73997
rect -1260 64140 42053 71660
rect 675498 70140 718860 154904
rect -1260 61660 41260 64140
rect 675547 63340 718860 70140
rect -1260 54140 42053 61660
rect 676340 60860 718860 63340
rect -1260 51660 40853 54140
rect 675547 53340 718860 60860
rect -1261 49277 41260 51660
rect -1261 40853 41560 49277
rect 43501 40853 63260 42960
rect 64881 41260 86283 42170
rect 109881 41260 131283 42170
rect 132881 41260 154283 42170
rect 155881 41260 177283 42170
rect 178881 41260 200283 42170
rect 204740 41260 212260 42053
rect 214740 41260 222260 42053
rect 64881 40853 86403 41260
rect 90616 40853 108363 41260
rect 109881 40853 131403 41260
rect 132881 40853 154403 41260
rect 155881 40853 177403 41260
rect 178881 40853 200403 41260
rect 204740 40853 222260 41260
rect 224501 40853 244260 42960
rect 248740 40860 266260 41660
rect 270740 40860 288260 41660
rect 292740 40860 310260 41660
rect 314740 40860 332260 41660
rect 336740 41260 344260 42053
rect 346740 41260 354260 42053
rect 248660 40853 266340 40860
rect 270660 40853 288340 40860
rect 292660 40853 310340 40860
rect 314660 40853 332340 40860
rect 336740 40853 354260 41260
rect 360501 40853 380260 42960
rect 381881 41260 403283 42170
rect 404881 41260 426283 42170
rect 427881 41260 449283 42170
rect 450881 41260 472283 42170
rect 476740 41260 484260 42053
rect 486740 41260 494260 42053
rect 381881 40853 403403 41260
rect 404881 40853 426403 41260
rect 427881 40853 449403 41260
rect 450881 40853 472403 41260
rect 476740 40853 494260 41260
rect 498740 41260 506260 42053
rect 508740 41260 516260 42053
rect 524740 41260 532260 42053
rect 534740 41260 542260 42053
rect 498740 40853 542260 41260
rect 548501 40853 568260 42960
rect 572740 40853 671260 52003
rect 676747 50860 718860 53340
rect 676340 49555 718861 50860
rect 676040 41260 718861 49555
rect 675540 40853 718861 41260
rect -1261 39540 718861 40853
rect -1260 38740 718861 39540
rect -1260 -1260 718860 38740
rect 572740 -1464 671260 -1260
<< metal1 >>
rect 101959 40130 101969 40330
rect 102023 40130 102033 40330
rect 101973 39934 102019 40130
<< via1 >>
rect 101969 40130 102023 40330
<< metal2 >>
rect 336566 997588 338362 997600
rect 336566 997212 336578 997588
rect 338350 997212 338362 997588
rect 67878 996690 68002 996890
rect 68468 996690 68520 996890
rect 68782 996690 68834 996890
rect 69102 996690 69154 996890
rect 70350 996690 70402 996890
rect 71061 996690 71113 996890
rect 72270 996690 72322 996890
rect 73119 996690 73171 996890
rect 73497 996690 73549 996890
rect 73848 996690 73900 996890
rect 74162 996690 74214 996890
rect 74891 996690 74943 996890
rect 75473 996690 75529 996890
rect 76848 996690 76900 996890
rect 77144 996690 77196 996890
rect 77770 996690 77822 996890
rect 80058 996690 80110 996890
rect 80362 996690 80576 996890
rect 81166 996690 81218 996890
rect 81454 996690 81584 996890
rect 82714 996690 82842 996890
rect 83090 996690 83142 996890
rect 83390 996690 83442 996890
rect 83688 996690 83740 996890
rect 83990 996690 84042 996890
rect 84290 996690 84342 996890
rect 85254 996690 85306 996890
rect 85616 996690 85668 996890
rect 91878 996690 92002 996890
rect 92468 996690 92520 996890
rect 92782 996690 92834 996890
rect 93102 996690 93154 996890
rect 94350 996690 94402 996890
rect 95061 996690 95113 996890
rect 96270 996690 96322 996890
rect 97119 996690 97171 996890
rect 97497 996690 97549 996890
rect 97848 996690 97900 996890
rect 98162 996690 98214 996890
rect 98891 996690 98943 996890
rect 99473 996690 99529 996890
rect 100848 996690 100900 996890
rect 101144 996690 101196 996890
rect 101770 996690 101822 996890
rect 104058 996690 104110 996890
rect 104362 996690 104576 996890
rect 105166 996690 105218 996890
rect 105454 996690 105584 996890
rect 106714 996690 106842 996890
rect 107090 996690 107142 996890
rect 107390 996690 107442 996890
rect 107688 996690 107740 996890
rect 107990 996690 108042 996890
rect 108290 996690 108342 996890
rect 109254 996690 109306 996890
rect 109616 996690 109668 996890
rect 115878 996690 116002 996890
rect 116468 996690 116520 996890
rect 116782 996690 116834 996890
rect 117102 996690 117154 996890
rect 118350 996690 118402 996890
rect 119061 996690 119113 996890
rect 120270 996690 120322 996890
rect 121119 996690 121171 996890
rect 121497 996690 121549 996890
rect 121848 996690 121900 996890
rect 122162 996690 122214 996890
rect 122891 996690 122943 996890
rect 123473 996690 123529 996890
rect 124848 996690 124900 996890
rect 125144 996690 125196 996890
rect 125770 996690 125822 996890
rect 128058 996690 128110 996890
rect 128362 996690 128576 996890
rect 129166 996690 129218 996890
rect 129454 996690 129584 996890
rect 130714 996690 130842 996890
rect 131090 996690 131142 996890
rect 131390 996690 131442 996890
rect 131688 996690 131740 996890
rect 131990 996690 132042 996890
rect 132290 996690 132342 996890
rect 133254 996690 133306 996890
rect 133616 996690 133668 996890
rect 139878 996690 140002 996890
rect 140468 996690 140520 996890
rect 140782 996690 140834 996890
rect 141102 996690 141154 996890
rect 142350 996690 142402 996890
rect 143061 996690 143113 996890
rect 144270 996690 144322 996890
rect 145119 996690 145171 996890
rect 145497 996690 145549 996890
rect 145848 996690 145900 996890
rect 146162 996690 146214 996890
rect 146891 996690 146943 996890
rect 147473 996690 147529 996890
rect 148848 996690 148900 996890
rect 149144 996690 149196 996890
rect 149770 996690 149822 996890
rect 152058 996690 152110 996890
rect 152362 996690 152576 996890
rect 153166 996690 153218 996890
rect 153454 996690 153584 996890
rect 154714 996690 154842 996890
rect 155090 996690 155142 996890
rect 155390 996690 155442 996890
rect 155688 996690 155740 996890
rect 155990 996690 156042 996890
rect 156290 996690 156342 996890
rect 157254 996690 157306 996890
rect 157616 996690 157668 996890
rect 209878 996690 210002 996890
rect 210468 996690 210520 996890
rect 210782 996690 210834 996890
rect 211102 996690 211154 996890
rect 212350 996690 212402 996890
rect 213061 996690 213113 996890
rect 214270 996690 214322 996890
rect 215119 996690 215171 996890
rect 215497 996690 215549 996890
rect 215848 996690 215900 996890
rect 216162 996690 216214 996890
rect 216891 996690 216943 996890
rect 217473 996690 217529 996890
rect 218848 996690 218900 996890
rect 219144 996690 219196 996890
rect 219770 996690 219822 996890
rect 222058 996690 222110 996890
rect 222362 996690 222576 996890
rect 223166 996690 223218 996890
rect 223454 996690 223584 996890
rect 224714 996690 224842 996890
rect 225090 996690 225142 996890
rect 225390 996690 225442 996890
rect 225688 996690 225740 996890
rect 225990 996690 226042 996890
rect 226290 996690 226342 996890
rect 227254 996690 227306 996890
rect 227616 996690 227668 996890
rect 233878 996690 234002 996890
rect 234468 996690 234520 996890
rect 234782 996690 234834 996890
rect 235102 996690 235154 996890
rect 236350 996690 236402 996890
rect 237061 996690 237113 996890
rect 238270 996690 238322 996890
rect 239119 996690 239171 996890
rect 239497 996690 239549 996890
rect 239848 996690 239900 996890
rect 240162 996690 240214 996890
rect 240891 996690 240943 996890
rect 241473 996690 241529 996890
rect 242848 996690 242900 996890
rect 243144 996690 243196 996890
rect 243770 996690 243822 996890
rect 246058 996690 246110 996890
rect 246362 996690 246576 996890
rect 247166 996690 247218 996890
rect 247454 996690 247584 996890
rect 248714 996690 248842 996890
rect 249090 996690 249142 996890
rect 249390 996690 249442 996890
rect 249688 996690 249740 996890
rect 249990 996690 250042 996890
rect 250290 996690 250342 996890
rect 251254 996690 251306 996890
rect 251616 996690 251668 996890
rect 257878 996690 258002 996890
rect 258468 996690 258520 996890
rect 258782 996690 258834 996890
rect 259102 996690 259154 996890
rect 260350 996690 260402 996890
rect 261061 996690 261113 996890
rect 262270 996690 262322 996890
rect 263119 996690 263171 996890
rect 263497 996690 263549 996890
rect 263848 996690 263900 996890
rect 264162 996690 264214 996890
rect 264891 996690 264943 996890
rect 265473 996690 265529 996890
rect 266848 996690 266900 996890
rect 267144 996690 267196 996890
rect 267770 996690 267822 996890
rect 270058 996690 270110 996890
rect 270362 996690 270576 996890
rect 271166 996690 271218 996890
rect 271454 996690 271584 996890
rect 272714 996690 272842 996890
rect 273090 996690 273142 996890
rect 273390 996690 273442 996890
rect 273688 996690 273740 996890
rect 273990 996690 274042 996890
rect 274290 996690 274342 996890
rect 275254 996690 275306 996890
rect 275616 996690 275668 996890
rect 281878 996690 282002 996890
rect 282468 996690 282520 996890
rect 282782 996690 282834 996890
rect 283102 996690 283154 996890
rect 284350 996690 284402 996890
rect 285061 996690 285113 996890
rect 286270 996690 286322 996890
rect 287119 996690 287171 996890
rect 287497 996690 287549 996890
rect 287848 996690 287900 996890
rect 288162 996690 288214 996890
rect 288891 996690 288943 996890
rect 289473 996690 289529 996890
rect 290848 996690 290900 996890
rect 291144 996690 291196 996890
rect 291770 996690 291822 996890
rect 294058 996690 294110 996890
rect 294362 996690 294576 996890
rect 295166 996690 295218 996890
rect 295454 996690 295584 996890
rect 296714 996690 296842 996890
rect 297090 996690 297142 996890
rect 297390 996690 297442 996890
rect 297688 996690 297740 996890
rect 297990 996690 298042 996890
rect 298290 996690 298342 996890
rect 299254 996690 299306 996890
rect 299616 996690 299668 996890
rect 336566 996600 338362 997212
rect 359566 997588 361362 997600
rect 359566 997212 359578 997588
rect 361350 997212 361362 997588
rect 359566 996600 361362 997212
rect 368496 996600 368624 997200
rect 368752 996600 368880 997200
rect 420878 996690 421002 996890
rect 421468 996690 421520 996890
rect 421782 996690 421834 996890
rect 422102 996690 422154 996890
rect 423350 996690 423402 996890
rect 424061 996690 424113 996890
rect 425270 996690 425322 996890
rect 426119 996690 426171 996890
rect 426497 996690 426549 996890
rect 426848 996690 426900 996890
rect 427162 996690 427214 996890
rect 427891 996690 427943 996890
rect 428473 996690 428529 996890
rect 429848 996690 429900 996890
rect 430144 996690 430196 996890
rect 430770 996690 430822 996890
rect 433058 996690 433110 996890
rect 433362 996690 433576 996890
rect 434166 996690 434218 996890
rect 434454 996690 434584 996890
rect 435714 996690 435842 996890
rect 436090 996690 436142 996890
rect 436390 996690 436442 996890
rect 436688 996690 436740 996890
rect 436990 996690 437042 996890
rect 437290 996690 437342 996890
rect 438254 996690 438306 996890
rect 438616 996690 438668 996890
rect 444878 996690 445002 996890
rect 445468 996690 445520 996890
rect 445782 996690 445834 996890
rect 446102 996690 446154 996890
rect 447350 996690 447402 996890
rect 448061 996690 448113 996890
rect 449270 996690 449322 996890
rect 450119 996690 450171 996890
rect 450497 996690 450549 996890
rect 450848 996690 450900 996890
rect 451162 996690 451214 996890
rect 451891 996690 451943 996890
rect 452473 996690 452529 996890
rect 453848 996690 453900 996890
rect 454144 996690 454196 996890
rect 454770 996690 454822 996890
rect 457058 996690 457110 996890
rect 457362 996690 457576 996890
rect 458166 996690 458218 996890
rect 458454 996690 458584 996890
rect 459714 996690 459842 996890
rect 460090 996690 460142 996890
rect 460390 996690 460442 996890
rect 460688 996690 460740 996890
rect 460990 996690 461042 996890
rect 461290 996690 461342 996890
rect 462254 996690 462306 996890
rect 462616 996690 462668 996890
rect 468878 996690 469002 996890
rect 469468 996690 469520 996890
rect 469782 996690 469834 996890
rect 470102 996690 470154 996890
rect 471350 996690 471402 996890
rect 472061 996690 472113 996890
rect 473270 996690 473322 996890
rect 474119 996690 474171 996890
rect 474497 996690 474549 996890
rect 474848 996690 474900 996890
rect 475162 996690 475214 996890
rect 475891 996690 475943 996890
rect 476473 996690 476529 996890
rect 477848 996690 477900 996890
rect 478144 996690 478196 996890
rect 478770 996690 478822 996890
rect 481058 996690 481110 996890
rect 481362 996690 481576 996890
rect 482166 996690 482218 996890
rect 482454 996690 482584 996890
rect 483714 996690 483842 996890
rect 484090 996690 484142 996890
rect 484390 996690 484442 996890
rect 484688 996690 484740 996890
rect 484990 996690 485042 996890
rect 485290 996690 485342 996890
rect 486254 996690 486306 996890
rect 486616 996690 486668 996890
rect 492878 996690 493002 996890
rect 493468 996690 493520 996890
rect 493782 996690 493834 996890
rect 494102 996690 494154 996890
rect 495350 996690 495402 996890
rect 496061 996690 496113 996890
rect 497270 996690 497322 996890
rect 498119 996690 498171 996890
rect 498497 996690 498549 996890
rect 498848 996690 498900 996890
rect 499162 996690 499214 996890
rect 499891 996690 499943 996890
rect 500473 996690 500529 996890
rect 501848 996690 501900 996890
rect 502144 996690 502196 996890
rect 502770 996690 502822 996890
rect 505058 996690 505110 996890
rect 505362 996690 505576 996890
rect 506166 996690 506218 996890
rect 506454 996690 506584 996890
rect 507714 996690 507842 996890
rect 508090 996690 508142 996890
rect 508390 996690 508442 996890
rect 508688 996690 508740 996890
rect 508990 996690 509042 996890
rect 509290 996690 509342 996890
rect 510254 996690 510306 996890
rect 510616 996690 510668 996890
rect 562878 996690 563002 996890
rect 563468 996690 563520 996890
rect 563782 996690 563834 996890
rect 564102 996690 564154 996890
rect 565350 996690 565402 996890
rect 566061 996690 566113 996890
rect 567270 996690 567322 996890
rect 568119 996690 568171 996890
rect 568497 996690 568549 996890
rect 568848 996690 568900 996890
rect 569162 996690 569214 996890
rect 569891 996690 569943 996890
rect 570473 996690 570529 996890
rect 571848 996690 571900 996890
rect 572144 996690 572196 996890
rect 572770 996690 572822 996890
rect 575058 996690 575110 996890
rect 575362 996690 575576 996890
rect 576166 996690 576218 996890
rect 576454 996690 576584 996890
rect 577714 996690 577842 996890
rect 578090 996690 578142 996890
rect 578390 996690 578442 996890
rect 578688 996690 578740 996890
rect 578990 996690 579042 996890
rect 579290 996690 579342 996890
rect 580254 996690 580306 996890
rect 580616 996690 580668 996890
rect 586878 996690 587002 996890
rect 587468 996690 587520 996890
rect 587782 996690 587834 996890
rect 588102 996690 588154 996890
rect 589350 996690 589402 996890
rect 590061 996690 590113 996890
rect 591270 996690 591322 996890
rect 592119 996690 592171 996890
rect 592497 996690 592549 996890
rect 592848 996690 592900 996890
rect 593162 996690 593214 996890
rect 593891 996690 593943 996890
rect 594473 996690 594529 996890
rect 595848 996690 595900 996890
rect 596144 996690 596196 996890
rect 596770 996690 596822 996890
rect 599058 996690 599110 996890
rect 599362 996690 599576 996890
rect 600166 996690 600218 996890
rect 600454 996690 600584 996890
rect 601714 996690 601842 996890
rect 602090 996690 602142 996890
rect 602390 996690 602442 996890
rect 602688 996690 602740 996890
rect 602990 996690 603042 996890
rect 603290 996690 603342 996890
rect 604254 996690 604306 996890
rect 604616 996690 604668 996890
rect 610878 996690 611002 996890
rect 611468 996690 611520 996890
rect 611782 996690 611834 996890
rect 612102 996690 612154 996890
rect 613350 996690 613402 996890
rect 614061 996690 614113 996890
rect 615270 996690 615322 996890
rect 616119 996690 616171 996890
rect 616497 996690 616549 996890
rect 616848 996690 616900 996890
rect 617162 996690 617214 996890
rect 617891 996690 617943 996890
rect 618473 996690 618529 996890
rect 619848 996690 619900 996890
rect 620144 996690 620196 996890
rect 620770 996690 620822 996890
rect 623058 996690 623110 996890
rect 623362 996690 623576 996890
rect 624166 996690 624218 996890
rect 624454 996690 624584 996890
rect 625714 996690 625842 996890
rect 626090 996690 626142 996890
rect 626390 996690 626442 996890
rect 626688 996690 626740 996890
rect 626990 996690 627042 996890
rect 627290 996690 627342 996890
rect 628254 996690 628306 996890
rect 628616 996690 628668 996890
rect 634878 996690 635002 996890
rect 635468 996690 635520 996890
rect 635782 996690 635834 996890
rect 636102 996690 636154 996890
rect 637350 996690 637402 996890
rect 638061 996690 638113 996890
rect 639270 996690 639322 996890
rect 640119 996690 640171 996890
rect 640497 996690 640549 996890
rect 640848 996690 640900 996890
rect 641162 996690 641214 996890
rect 641891 996690 641943 996890
rect 642473 996690 642529 996890
rect 643848 996690 643900 996890
rect 644144 996690 644196 996890
rect 644770 996690 644822 996890
rect 647058 996690 647110 996890
rect 647362 996690 647576 996890
rect 648166 996690 648218 996890
rect 648454 996690 648584 996890
rect 649714 996690 649842 996890
rect 650090 996690 650142 996890
rect 650390 996690 650442 996890
rect 650688 996690 650740 996890
rect 650990 996690 651042 996890
rect 651290 996690 651342 996890
rect 652254 996690 652306 996890
rect 652616 996690 652668 996890
rect 576666 50743 576794 51343
rect 576966 50743 577094 51343
rect 579167 50743 579219 51343
rect 579317 50743 579369 51343
rect 579467 50743 579519 51343
rect 579617 50743 579669 51343
rect 579772 50743 579814 51343
rect 579926 50743 579962 51343
rect 580073 50743 580116 51343
rect 580217 50743 580269 51343
rect 580367 50743 580419 51343
rect 580980 50743 581032 51343
rect 585410 50743 585462 51343
rect 586059 50743 586111 51343
rect 588949 50743 589001 51343
rect 589380 50743 589432 51343
rect 609051 50743 609220 51343
rect 609249 50743 609418 51343
rect 613341 50743 613393 51343
rect 614017 50743 614069 51343
rect 616290 50743 616342 51343
rect 617624 50743 617676 51343
rect 619034 50743 619086 51343
rect 619114 50743 619166 51343
rect 620239 50743 620308 51343
rect 620400 50743 620452 51343
rect 620480 50743 620532 51343
rect 621442 50743 621494 51343
rect 621522 50743 621574 51343
rect 621960 50743 622012 51343
rect 622681 50743 622733 51343
rect 622761 50743 622813 51343
rect 623195 50743 623247 51343
rect 623275 50743 623327 51343
rect 627397 50743 627797 51343
rect 634202 50743 634602 51343
rect 638672 50743 638724 51343
rect 638752 50743 638804 51343
rect 639186 50743 639238 51343
rect 639987 50743 640039 51343
rect 640425 50743 640477 51343
rect 640505 50743 640557 51343
rect 641467 50743 641519 51343
rect 641547 50743 641599 51343
rect 641691 50743 641760 51343
rect 642833 50743 642885 51343
rect 642913 50743 642965 51343
rect 644323 50743 644375 51343
rect 645657 50743 645709 51343
rect 647930 50743 647982 51343
rect 648606 50743 648658 51343
rect 652581 50743 652751 51343
rect 652779 50743 652948 51343
rect 67131 40710 67183 40910
rect 67493 40710 67545 40910
rect 68457 40710 68509 40910
rect 68757 40710 68809 40910
rect 69059 40710 69111 40910
rect 69357 40710 69409 40910
rect 69657 40710 69709 40910
rect 69957 40710 70085 40910
rect 71215 40710 71345 40910
rect 71581 40710 71633 40910
rect 72223 40710 72437 40910
rect 72689 40710 72741 40910
rect 74977 40710 75029 40910
rect 75603 40710 75655 40910
rect 75899 40710 75951 40910
rect 77270 40710 77326 40910
rect 77856 40710 77908 40910
rect 78585 40710 78637 40910
rect 78899 40710 78951 40910
rect 79250 40710 79302 40910
rect 79628 40710 79680 40910
rect 80477 40710 80529 40910
rect 81686 40710 81738 40910
rect 82397 40710 82449 40910
rect 83645 40710 83697 40910
rect 83965 40710 84017 40910
rect 84279 40710 84331 40910
rect 84797 40710 84921 40910
rect 112131 40710 112183 40910
rect 112493 40710 112545 40910
rect 113457 40710 113509 40910
rect 113757 40710 113809 40910
rect 114059 40710 114111 40910
rect 114357 40710 114409 40910
rect 114657 40710 114709 40910
rect 114957 40710 115085 40910
rect 116215 40710 116345 40910
rect 116581 40710 116633 40910
rect 117223 40710 117437 40910
rect 117689 40710 117741 40910
rect 119977 40710 120029 40910
rect 120603 40710 120655 40910
rect 120899 40710 120951 40910
rect 122270 40710 122326 40910
rect 122856 40710 122908 40910
rect 123585 40710 123637 40910
rect 123899 40710 123951 40910
rect 124250 40710 124302 40910
rect 124628 40710 124680 40910
rect 125477 40710 125529 40910
rect 126686 40710 126738 40910
rect 127397 40710 127449 40910
rect 128645 40710 128697 40910
rect 128965 40710 129017 40910
rect 129279 40710 129331 40910
rect 129797 40710 129921 40910
rect 135131 40710 135183 40910
rect 135493 40710 135545 40910
rect 136457 40710 136509 40910
rect 136757 40710 136809 40910
rect 137059 40710 137111 40910
rect 137357 40710 137409 40910
rect 137657 40710 137709 40910
rect 137957 40710 138085 40910
rect 139215 40710 139345 40910
rect 139581 40710 139633 40910
rect 140223 40710 140437 40910
rect 140689 40710 140741 40910
rect 142977 40710 143029 40910
rect 143603 40710 143655 40910
rect 143899 40710 143951 40910
rect 145270 40710 145326 40910
rect 145856 40710 145908 40910
rect 146585 40710 146637 40910
rect 146899 40710 146951 40910
rect 147250 40710 147302 40910
rect 147628 40710 147680 40910
rect 148477 40710 148529 40910
rect 149686 40710 149738 40910
rect 150397 40710 150449 40910
rect 151645 40710 151697 40910
rect 151965 40710 152017 40910
rect 152279 40710 152331 40910
rect 152797 40710 152921 40910
rect 158131 40710 158183 40910
rect 158493 40710 158545 40910
rect 159457 40710 159509 40910
rect 159757 40710 159809 40910
rect 160059 40710 160111 40910
rect 160357 40710 160409 40910
rect 160657 40710 160709 40910
rect 160957 40710 161085 40910
rect 162215 40710 162345 40910
rect 162581 40710 162633 40910
rect 163223 40710 163437 40910
rect 163689 40710 163741 40910
rect 165977 40710 166029 40910
rect 166603 40710 166655 40910
rect 166899 40710 166951 40910
rect 168270 40710 168326 40910
rect 168856 40710 168908 40910
rect 169585 40710 169637 40910
rect 169899 40710 169951 40910
rect 170250 40710 170302 40910
rect 170628 40710 170680 40910
rect 171477 40710 171529 40910
rect 172686 40710 172738 40910
rect 173397 40710 173449 40910
rect 174645 40710 174697 40910
rect 174965 40710 175017 40910
rect 175279 40710 175331 40910
rect 175797 40710 175921 40910
rect 181131 40710 181183 40910
rect 181493 40710 181545 40910
rect 182457 40710 182509 40910
rect 182757 40710 182809 40910
rect 183059 40710 183111 40910
rect 183357 40710 183409 40910
rect 183657 40710 183709 40910
rect 183957 40710 184085 40910
rect 185215 40710 185345 40910
rect 185581 40710 185633 40910
rect 186223 40710 186437 40910
rect 186689 40710 186741 40910
rect 188977 40710 189029 40910
rect 189603 40710 189655 40910
rect 189899 40710 189951 40910
rect 191270 40710 191326 40910
rect 191856 40710 191908 40910
rect 192585 40710 192637 40910
rect 192899 40710 192951 40910
rect 193250 40710 193302 40910
rect 193628 40710 193680 40910
rect 194477 40710 194529 40910
rect 195686 40710 195738 40910
rect 196397 40710 196449 40910
rect 197645 40710 197697 40910
rect 197965 40710 198017 40910
rect 198279 40710 198331 40910
rect 198797 40710 198921 40910
rect 92353 40000 92557 40600
rect 100396 40000 100448 40600
rect 100769 40000 100899 40600
rect 101067 40000 101213 40600
rect 101354 40000 101484 40600
rect 101969 40330 102023 40600
rect 101969 40120 102023 40130
rect 102468 40000 102528 40600
rect 102755 40000 102985 40600
rect 103218 40000 103551 40600
rect 103973 40000 104089 40600
rect 104491 40000 104543 40600
rect 105221 40000 105315 40600
rect 255438 40388 257234 41000
rect 255438 40012 255450 40388
rect 257222 40012 257234 40388
rect 255438 40000 257234 40012
rect 277438 40388 279234 41000
rect 277438 40012 277450 40388
rect 279222 40012 279234 40388
rect 277438 40000 279234 40012
rect 299438 40388 301234 41000
rect 299438 40012 299450 40388
rect 301222 40012 301234 40388
rect 299438 40000 301234 40012
rect 321438 40388 323234 41000
rect 384131 40710 384183 40910
rect 384493 40710 384545 40910
rect 385457 40710 385509 40910
rect 385757 40710 385809 40910
rect 386059 40710 386111 40910
rect 386357 40710 386409 40910
rect 386657 40710 386709 40910
rect 386957 40710 387085 40910
rect 388215 40710 388345 40910
rect 388581 40710 388633 40910
rect 389223 40710 389437 40910
rect 389689 40710 389741 40910
rect 391977 40710 392029 40910
rect 392603 40710 392655 40910
rect 392899 40710 392951 40910
rect 394270 40710 394326 40910
rect 394856 40710 394908 40910
rect 395585 40710 395637 40910
rect 395899 40710 395951 40910
rect 396250 40710 396302 40910
rect 396628 40710 396680 40910
rect 397477 40710 397529 40910
rect 398686 40710 398738 40910
rect 399397 40710 399449 40910
rect 400645 40710 400697 40910
rect 400965 40710 401017 40910
rect 401279 40710 401331 40910
rect 401797 40710 401921 40910
rect 407131 40710 407183 40910
rect 407493 40710 407545 40910
rect 408457 40710 408509 40910
rect 408757 40710 408809 40910
rect 409059 40710 409111 40910
rect 409357 40710 409409 40910
rect 409657 40710 409709 40910
rect 409957 40710 410085 40910
rect 411215 40710 411345 40910
rect 411581 40710 411633 40910
rect 412223 40710 412437 40910
rect 412689 40710 412741 40910
rect 414977 40710 415029 40910
rect 415603 40710 415655 40910
rect 415899 40710 415951 40910
rect 417270 40710 417326 40910
rect 417856 40710 417908 40910
rect 418585 40710 418637 40910
rect 418899 40710 418951 40910
rect 419250 40710 419302 40910
rect 419628 40710 419680 40910
rect 420477 40710 420529 40910
rect 421686 40710 421738 40910
rect 422397 40710 422449 40910
rect 423645 40710 423697 40910
rect 423965 40710 424017 40910
rect 424279 40710 424331 40910
rect 424797 40710 424921 40910
rect 430131 40710 430183 40910
rect 430493 40710 430545 40910
rect 431457 40710 431509 40910
rect 431757 40710 431809 40910
rect 432059 40710 432111 40910
rect 432357 40710 432409 40910
rect 432657 40710 432709 40910
rect 432957 40710 433085 40910
rect 434215 40710 434345 40910
rect 434581 40710 434633 40910
rect 435223 40710 435437 40910
rect 435689 40710 435741 40910
rect 437977 40710 438029 40910
rect 438603 40710 438655 40910
rect 438899 40710 438951 40910
rect 440270 40710 440326 40910
rect 440856 40710 440908 40910
rect 441585 40710 441637 40910
rect 441899 40710 441951 40910
rect 442250 40710 442302 40910
rect 442628 40710 442680 40910
rect 443477 40710 443529 40910
rect 444686 40710 444738 40910
rect 445397 40710 445449 40910
rect 446645 40710 446697 40910
rect 446965 40710 447017 40910
rect 447279 40710 447331 40910
rect 447797 40710 447921 40910
rect 453131 40710 453183 40910
rect 453493 40710 453545 40910
rect 454457 40710 454509 40910
rect 454757 40710 454809 40910
rect 455059 40710 455111 40910
rect 455357 40710 455409 40910
rect 455657 40710 455709 40910
rect 455957 40710 456085 40910
rect 457215 40710 457345 40910
rect 457581 40710 457633 40910
rect 458223 40710 458437 40910
rect 458689 40710 458741 40910
rect 460977 40710 461029 40910
rect 461603 40710 461655 40910
rect 461899 40710 461951 40910
rect 463270 40710 463326 40910
rect 463856 40710 463908 40910
rect 464585 40710 464637 40910
rect 464899 40710 464951 40910
rect 465250 40710 465302 40910
rect 465628 40710 465680 40910
rect 466477 40710 466529 40910
rect 467686 40710 467738 40910
rect 468397 40710 468449 40910
rect 469645 40710 469697 40910
rect 469965 40710 470017 40910
rect 470279 40710 470331 40910
rect 470797 40710 470921 40910
rect 321438 40012 321450 40388
rect 323222 40012 323234 40388
rect 321438 40000 323234 40012
rect 515865 40000 515917 40600
rect 516097 40000 516149 40600
rect 516344 40000 516396 40600
rect 516556 40000 516608 40600
rect 516896 40000 516948 40600
rect 517210 40000 517262 40600
rect 517427 40000 517479 40600
rect 517659 40000 517711 40600
rect 517952 40000 518004 40600
rect 519285 40000 519337 40600
rect 523619 40000 523697 40600
rect 523965 40000 524017 40600
rect 524219 40000 524271 40600
rect 524476 40000 524528 40600
rect 524713 40000 524765 40600
rect 525846 40000 525898 40600
<< via2 >>
rect 336578 997212 338350 997588
rect 359578 997212 361350 997588
rect 255450 40012 257222 40388
rect 277450 40012 279222 40388
rect 299450 40012 301222 40388
rect 321450 40012 323222 40388
<< metal3 >>
rect 44898 996807 49700 998007
rect 49990 996807 54652 997807
rect 54951 996807 59740 998007
rect 163899 996807 168679 998007
rect 173878 996807 178658 998007
rect 186900 996807 191700 998007
rect 192000 997807 194176 998007
rect 194476 997807 196651 998007
rect 192000 996807 196651 997807
rect 196951 996807 201740 998007
rect 305899 996807 310679 998007
rect 315878 996807 320658 998007
rect 336566 997588 338362 998000
rect 336566 997212 336578 997588
rect 338350 997212 338362 997588
rect 336566 997200 338362 997212
rect 359566 997588 361362 998000
rect 359566 997212 359578 997588
rect 361350 997212 361362 997588
rect 359566 997200 361362 997212
rect 374899 996807 379679 998007
rect 384878 996807 389658 998007
rect 397899 996807 402679 998007
rect 407878 996807 412658 998007
rect 516898 996807 521700 998007
rect 521990 996807 526652 997807
rect 526951 996807 531740 998007
rect 539899 996807 544679 998007
rect 549878 996807 554658 998007
rect 658900 996807 663700 998007
rect 664000 997807 666176 998007
rect 666476 997807 668651 998007
rect 664000 996807 668651 997807
rect 668951 996807 673740 998007
rect 676700 995432 677300 995492
rect 40300 995154 40900 995214
rect 676700 995096 677300 995156
rect 676700 994844 677300 994904
rect 676700 994592 677300 994652
rect 676700 994340 677300 994400
rect 40300 994274 40900 994334
rect 676700 994088 677300 994148
rect 40300 990652 40900 990712
rect 676700 990466 677300 990526
rect 40300 990400 40900 990460
rect 40300 990148 40900 990208
rect 40300 989896 40900 989956
rect 40300 989644 40900 989704
rect 676700 989586 677300 989646
rect 40300 989308 40900 989368
rect 39593 982078 40793 986858
rect 676807 981321 678007 986101
rect 39593 972099 40793 976879
rect 676807 971342 678007 976122
rect 39593 959151 40793 963940
rect 39593 956676 40793 958851
rect 676807 957300 678007 962102
rect 39793 956376 40793 956676
rect 39593 954200 40793 956376
rect 39593 949100 40793 953900
rect 676807 952348 677807 957010
rect 676807 947260 678007 952049
rect 40542 946252 40842 946322
rect 40542 945802 40842 945872
rect 40542 944602 40842 944672
rect 40542 944304 40842 944374
rect 40538 944024 40838 944094
rect 40542 943712 40842 943782
rect 40542 943438 40842 943508
rect 40542 943090 40842 943218
rect 676758 941996 677058 942120
rect 40542 941658 40842 941788
rect 676758 941468 677058 941538
rect 40542 941128 40842 941198
rect 676758 941058 677058 941128
rect 40542 940564 40842 940778
rect 676758 940714 677058 940784
rect 40542 939932 40842 940002
rect 676758 939852 677058 939922
rect 676758 939132 677058 939202
rect 676758 937932 677058 938002
rect 40542 937720 40842 937790
rect 40542 937172 40842 937242
rect 676758 937160 677058 937230
rect 676758 936676 677058 936746
rect 40542 936592 40842 936662
rect 676758 936232 677058 936302
rect 676758 935614 677058 935684
rect 40542 935426 40842 935496
rect 676758 935160 677058 935230
rect 40542 934970 40842 935040
rect 676758 934704 677058 934774
rect 40542 934516 40842 934586
rect 40542 933898 40842 933968
rect 676758 933538 677058 933608
rect 40542 933454 40842 933524
rect 40542 932970 40842 933040
rect 676758 932958 677058 933028
rect 676758 932410 677058 932480
rect 40542 932198 40842 932268
rect 40542 930998 40842 931068
rect 40542 930278 40842 930348
rect 676758 930198 677058 930268
rect 40542 929416 40842 929486
rect 676758 929422 677058 929636
rect 40542 929072 40842 929142
rect 676758 929002 677058 929072
rect 40542 928662 40842 928732
rect 676758 928412 677058 928542
rect 40542 928080 40842 928204
rect 676758 926982 677058 927110
rect 676758 926692 677058 926762
rect 676758 926418 677058 926488
rect 676762 926106 677062 926176
rect 676758 925826 677058 925896
rect 676758 925528 677058 925598
rect 40542 925252 40842 925322
rect 40542 924802 40842 924872
rect 676758 924328 677058 924398
rect 676758 923878 677058 923948
rect 40542 923602 40842 923672
rect 40542 923304 40842 923374
rect 40538 923024 40838 923094
rect 40542 922712 40842 922782
rect 40542 922438 40842 922508
rect 40542 922090 40842 922218
rect 676758 920996 677058 921120
rect 40542 920658 40842 920788
rect 676758 920468 677058 920538
rect 40542 920128 40842 920198
rect 676758 920058 677058 920128
rect 40542 919564 40842 919778
rect 676758 919714 677058 919784
rect 40542 918932 40842 919002
rect 676758 918852 677058 918922
rect 676758 918132 677058 918202
rect 676758 916932 677058 917002
rect 40542 916720 40842 916790
rect 40542 916172 40842 916242
rect 676758 916160 677058 916230
rect 676758 915676 677058 915746
rect 40542 915592 40842 915662
rect 676758 915232 677058 915302
rect 676758 914614 677058 914684
rect 40542 914426 40842 914496
rect 676758 914160 677058 914230
rect 40542 913970 40842 914040
rect 676758 913704 677058 913774
rect 40542 913516 40842 913586
rect 40542 912898 40842 912968
rect 676758 912538 677058 912608
rect 40542 912454 40842 912524
rect 40542 911970 40842 912040
rect 676758 911958 677058 912028
rect 676758 911410 677058 911480
rect 40542 911198 40842 911268
rect 40542 909998 40842 910068
rect 40542 909278 40842 909348
rect 676758 909198 677058 909268
rect 40542 908416 40842 908486
rect 676758 908422 677058 908636
rect 40542 908072 40842 908142
rect 676758 908002 677058 908072
rect 40542 907662 40842 907732
rect 676758 907412 677058 907542
rect 40542 907080 40842 907204
rect 676758 905982 677058 906110
rect 676758 905692 677058 905762
rect 676758 905418 677058 905488
rect 676762 905106 677062 905176
rect 676758 904826 677058 904896
rect 676758 904528 677058 904598
rect 40542 904252 40842 904322
rect 40542 903802 40842 903872
rect 676758 903328 677058 903398
rect 676758 902878 677058 902948
rect 40542 902602 40842 902672
rect 40542 902304 40842 902374
rect 40538 902024 40838 902094
rect 40542 901712 40842 901782
rect 40542 901438 40842 901508
rect 40542 901090 40842 901218
rect 676758 899996 677058 900120
rect 40542 899658 40842 899788
rect 676758 899468 677058 899538
rect 40542 899128 40842 899198
rect 676758 899058 677058 899128
rect 40542 898564 40842 898778
rect 676758 898714 677058 898784
rect 40542 897932 40842 898002
rect 676758 897852 677058 897922
rect 676758 897132 677058 897202
rect 676758 895932 677058 896002
rect 40542 895720 40842 895790
rect 40542 895172 40842 895242
rect 676758 895160 677058 895230
rect 676758 894676 677058 894746
rect 40542 894592 40842 894662
rect 676758 894232 677058 894302
rect 676758 893614 677058 893684
rect 40542 893426 40842 893496
rect 676758 893160 677058 893230
rect 40542 892970 40842 893040
rect 676758 892704 677058 892774
rect 40542 892516 40842 892586
rect 40542 891898 40842 891968
rect 676758 891538 677058 891608
rect 40542 891454 40842 891524
rect 40542 890970 40842 891040
rect 676758 890958 677058 891028
rect 676758 890410 677058 890480
rect 40542 890198 40842 890268
rect 40542 888998 40842 889068
rect 40542 888278 40842 888348
rect 676758 888198 677058 888268
rect 40542 887416 40842 887486
rect 676758 887422 677058 887636
rect 40542 887072 40842 887142
rect 676758 887002 677058 887072
rect 40542 886662 40842 886732
rect 676758 886412 677058 886542
rect 40542 886080 40842 886204
rect 676758 884982 677058 885110
rect 676758 884692 677058 884762
rect 676758 884418 677058 884488
rect 676762 884106 677062 884176
rect 676758 883826 677058 883896
rect 676758 883528 677058 883598
rect 40542 883252 40842 883322
rect 40542 882802 40842 882872
rect 676758 882328 677058 882398
rect 676758 881878 677058 881948
rect 40542 881602 40842 881672
rect 40542 881304 40842 881374
rect 40538 881024 40838 881094
rect 40542 880712 40842 880782
rect 40542 880438 40842 880508
rect 40542 880090 40842 880218
rect 676758 878996 677058 879120
rect 40542 878658 40842 878788
rect 676758 878468 677058 878538
rect 40542 878128 40842 878198
rect 676758 878058 677058 878128
rect 40542 877564 40842 877778
rect 676758 877714 677058 877784
rect 40542 876932 40842 877002
rect 676758 876852 677058 876922
rect 676758 876132 677058 876202
rect 676758 874932 677058 875002
rect 40542 874720 40842 874790
rect 40542 874172 40842 874242
rect 676758 874160 677058 874230
rect 676758 873676 677058 873746
rect 40542 873592 40842 873662
rect 676758 873232 677058 873302
rect 676758 872614 677058 872684
rect 40542 872426 40842 872496
rect 676758 872160 677058 872230
rect 40542 871970 40842 872040
rect 676758 871704 677058 871774
rect 40542 871516 40842 871586
rect 40542 870898 40842 870968
rect 676758 870538 677058 870608
rect 40542 870454 40842 870524
rect 40542 869970 40842 870040
rect 676758 869958 677058 870028
rect 676758 869410 677058 869480
rect 40542 869198 40842 869268
rect 40542 867998 40842 868068
rect 40542 867278 40842 867348
rect 676758 867198 677058 867268
rect 40542 866416 40842 866486
rect 676758 866422 677058 866636
rect 40542 866072 40842 866142
rect 676758 866002 677058 866072
rect 40542 865662 40842 865732
rect 676758 865412 677058 865542
rect 40542 865080 40842 865204
rect 676758 863982 677058 864110
rect 676758 863692 677058 863762
rect 676758 863418 677058 863488
rect 676762 863106 677062 863176
rect 676758 862826 677058 862896
rect 676758 862528 677058 862598
rect 676758 861328 677058 861398
rect 676758 860878 677058 860948
rect 39593 855078 40793 859858
rect 676807 853321 678007 858101
rect 39593 845099 40793 849879
rect 676807 843342 678007 848122
rect 40542 842252 40842 842322
rect 40542 841802 40842 841872
rect 40542 840602 40842 840672
rect 40542 840304 40842 840374
rect 40538 840024 40838 840094
rect 40542 839712 40842 839782
rect 40542 839438 40842 839508
rect 40542 839090 40842 839218
rect 676758 837996 677058 838120
rect 40542 837658 40842 837788
rect 676758 837468 677058 837538
rect 40542 837128 40842 837198
rect 676758 837058 677058 837128
rect 40542 836564 40842 836778
rect 676758 836714 677058 836784
rect 40542 835932 40842 836002
rect 676758 835852 677058 835922
rect 676758 835132 677058 835202
rect 676758 833932 677058 834002
rect 40542 833720 40842 833790
rect 40542 833172 40842 833242
rect 676758 833160 677058 833230
rect 676758 832676 677058 832746
rect 40542 832592 40842 832662
rect 676758 832232 677058 832302
rect 676758 831614 677058 831684
rect 40542 831426 40842 831496
rect 676758 831160 677058 831230
rect 40542 830970 40842 831040
rect 676758 830704 677058 830774
rect 40542 830516 40842 830586
rect 40542 829898 40842 829968
rect 676758 829538 677058 829608
rect 40542 829454 40842 829524
rect 40542 828970 40842 829040
rect 676758 828958 677058 829028
rect 676758 828410 677058 828480
rect 40542 828198 40842 828268
rect 40542 826998 40842 827068
rect 40542 826278 40842 826348
rect 676758 826198 677058 826268
rect 40542 825416 40842 825486
rect 676758 825422 677058 825636
rect 40542 825072 40842 825142
rect 676758 825002 677058 825072
rect 40542 824662 40842 824732
rect 676758 824412 677058 824542
rect 40542 824080 40842 824204
rect 676758 822982 677058 823110
rect 676758 822692 677058 822762
rect 676758 822418 677058 822488
rect 676762 822106 677062 822176
rect 676758 821826 677058 821896
rect 676758 821528 677058 821598
rect 40542 821252 40842 821322
rect 40542 820802 40842 820872
rect 676758 820328 677058 820398
rect 676758 819878 677058 819948
rect 40542 819602 40842 819672
rect 40542 819304 40842 819374
rect 40538 819024 40838 819094
rect 40542 818712 40842 818782
rect 40542 818438 40842 818508
rect 40542 818090 40842 818218
rect 676758 816996 677058 817120
rect 40542 816658 40842 816788
rect 676758 816468 677058 816538
rect 40542 816128 40842 816198
rect 676758 816058 677058 816128
rect 40542 815564 40842 815778
rect 676758 815714 677058 815784
rect 40542 814932 40842 815002
rect 676758 814852 677058 814922
rect 676758 814132 677058 814202
rect 676758 812932 677058 813002
rect 40542 812720 40842 812790
rect 40542 812172 40842 812242
rect 676758 812160 677058 812230
rect 676758 811676 677058 811746
rect 40542 811592 40842 811662
rect 676758 811232 677058 811302
rect 676758 810614 677058 810684
rect 40542 810426 40842 810496
rect 676758 810160 677058 810230
rect 40542 809970 40842 810040
rect 676758 809704 677058 809774
rect 40542 809516 40842 809586
rect 40542 808898 40842 808968
rect 676758 808538 677058 808608
rect 40542 808454 40842 808524
rect 40542 807970 40842 808040
rect 676758 807958 677058 808028
rect 676758 807410 677058 807480
rect 40542 807198 40842 807268
rect 40542 805998 40842 806068
rect 40542 805278 40842 805348
rect 676758 805198 677058 805268
rect 40542 804416 40842 804486
rect 676758 804422 677058 804636
rect 40542 804072 40842 804142
rect 676758 804002 677058 804072
rect 40542 803662 40842 803732
rect 676758 803412 677058 803542
rect 40542 803080 40842 803204
rect 676758 801982 677058 802110
rect 676758 801692 677058 801762
rect 676758 801418 677058 801488
rect 676762 801106 677062 801176
rect 676758 800826 677058 800896
rect 676758 800528 677058 800598
rect 40542 800252 40842 800322
rect 40542 799802 40842 799872
rect 676758 799328 677058 799398
rect 676758 798878 677058 798948
rect 40542 798602 40842 798672
rect 40542 798304 40842 798374
rect 40538 798024 40838 798094
rect 40542 797712 40842 797782
rect 40542 797438 40842 797508
rect 40542 797090 40842 797218
rect 676758 795996 677058 796120
rect 40542 795658 40842 795788
rect 676758 795468 677058 795538
rect 40542 795128 40842 795198
rect 676758 795058 677058 795128
rect 40542 794564 40842 794778
rect 676758 794714 677058 794784
rect 40542 793932 40842 794002
rect 676758 793852 677058 793922
rect 676758 793132 677058 793202
rect 676758 791932 677058 792002
rect 40542 791720 40842 791790
rect 40542 791172 40842 791242
rect 676758 791160 677058 791230
rect 676758 790676 677058 790746
rect 40542 790592 40842 790662
rect 676758 790232 677058 790302
rect 676758 789614 677058 789684
rect 40542 789426 40842 789496
rect 676758 789160 677058 789230
rect 40542 788970 40842 789040
rect 676758 788704 677058 788774
rect 40542 788516 40842 788586
rect 40542 787898 40842 787968
rect 676758 787538 677058 787608
rect 40542 787454 40842 787524
rect 40542 786970 40842 787040
rect 676758 786958 677058 787028
rect 676758 786410 677058 786480
rect 40542 786198 40842 786268
rect 40542 784998 40842 785068
rect 40542 784278 40842 784348
rect 676758 784198 677058 784268
rect 40542 783416 40842 783486
rect 676758 783422 677058 783636
rect 40542 783072 40842 783142
rect 676758 783002 677058 783072
rect 40542 782662 40842 782732
rect 676758 782412 677058 782542
rect 40542 782080 40842 782204
rect 676758 780982 677058 781110
rect 676758 780692 677058 780762
rect 676758 780418 677058 780488
rect 676762 780106 677062 780176
rect 676758 779826 677058 779896
rect 676758 779528 677058 779598
rect 40542 779252 40842 779322
rect 40542 778802 40842 778872
rect 676758 778328 677058 778398
rect 676758 777878 677058 777948
rect 40542 777602 40842 777672
rect 40542 777304 40842 777374
rect 40538 777024 40838 777094
rect 40542 776712 40842 776782
rect 40542 776438 40842 776508
rect 40542 776090 40842 776218
rect 676758 774996 677058 775120
rect 40542 774658 40842 774788
rect 676758 774468 677058 774538
rect 40542 774128 40842 774198
rect 676758 774058 677058 774128
rect 40542 773564 40842 773778
rect 676758 773714 677058 773784
rect 40542 772932 40842 773002
rect 676758 772852 677058 772922
rect 676758 772132 677058 772202
rect 676758 770932 677058 771002
rect 40542 770720 40842 770790
rect 40542 770172 40842 770242
rect 676758 770160 677058 770230
rect 676758 769676 677058 769746
rect 40542 769592 40842 769662
rect 676758 769232 677058 769302
rect 676758 768614 677058 768684
rect 40542 768426 40842 768496
rect 676758 768160 677058 768230
rect 40542 767970 40842 768040
rect 676758 767704 677058 767774
rect 40542 767516 40842 767586
rect 40542 766898 40842 766968
rect 676758 766538 677058 766608
rect 40542 766454 40842 766524
rect 40542 765970 40842 766040
rect 676758 765958 677058 766028
rect 676758 765410 677058 765480
rect 40542 765198 40842 765268
rect 40542 763998 40842 764068
rect 40542 763278 40842 763348
rect 676758 763198 677058 763268
rect 40542 762416 40842 762486
rect 676758 762422 677058 762636
rect 40542 762072 40842 762142
rect 676758 762002 677058 762072
rect 40542 761662 40842 761732
rect 676758 761412 677058 761542
rect 40542 761080 40842 761204
rect 676758 759982 677058 760110
rect 676758 759692 677058 759762
rect 676758 759418 677058 759488
rect 676762 759106 677062 759176
rect 676758 758826 677058 758896
rect 676758 758528 677058 758598
rect 676758 757328 677058 757398
rect 676758 756878 677058 756948
rect 39593 751151 40793 755940
rect 39793 746190 40793 750852
rect 676807 749300 678007 754100
rect 676807 746824 678007 749000
rect 676807 746524 677807 746824
rect 39593 741098 40793 745900
rect 676807 744349 678007 746524
rect 676807 739260 678007 744049
rect 39593 731078 40793 735858
rect 676807 729321 678007 734101
rect 39593 721099 40793 725879
rect 676807 719342 678007 724122
rect 39593 708078 40793 712858
rect 676807 705321 678007 710101
rect 39593 698099 40793 702879
rect 676807 695342 678007 700122
rect 39593 688078 40793 692858
rect 676807 685321 678007 690101
rect 39593 678099 40793 682879
rect 676807 675342 678007 680122
rect 40300 675252 40600 675322
rect 40300 674802 40600 674872
rect 40000 670995 40600 671061
rect 40000 670825 40600 670891
rect 40000 670655 40600 670721
rect 40000 670028 40600 670094
rect 677000 670014 677600 670134
rect 40000 669889 40600 669955
rect 677000 669760 677600 669879
rect 677000 669503 677600 669623
rect 677000 668927 677600 669047
rect 677000 668712 677600 668778
rect 677000 668511 677600 668577
rect 677000 668380 677600 668446
rect 40000 668058 40600 668178
rect 40000 666679 40600 666745
rect 40000 666509 40600 666575
rect 677000 666207 677600 666273
rect 677000 666058 677600 666124
rect 677000 665707 677600 665773
rect 677000 665258 677600 665324
rect 677000 664663 677600 664729
rect 40000 664169 40600 664243
rect 40000 662533 40600 662599
rect 40000 662363 40600 662429
rect 677000 661327 677600 661393
rect 677000 661063 677600 661129
rect 677000 660893 677600 660959
rect 40000 659825 40600 659891
rect 677000 659803 677600 659869
rect 40000 658387 40600 658453
rect 40000 658217 40600 658283
rect 40000 658047 40600 658113
rect 677000 657087 677600 657153
rect 677000 656917 677600 656983
rect 677000 656747 677600 656813
rect 40000 655331 40600 655397
rect 677000 655309 677600 655375
rect 40000 654241 40600 654307
rect 40000 654071 40600 654137
rect 40000 653807 40600 653873
rect 677000 652771 677600 652837
rect 677000 652601 677600 652667
rect 677000 650957 677600 651031
rect 40000 650471 40600 650537
rect 40000 649876 40600 649942
rect 40000 649427 40600 649493
rect 40000 649076 40600 649142
rect 40000 648927 40600 648993
rect 677000 648625 677600 648691
rect 677000 648455 677600 648521
rect 677000 647022 677600 647142
rect 40000 646754 40600 646820
rect 40000 646623 40600 646689
rect 40000 646422 40600 646488
rect 40000 646153 40600 646273
rect 40000 645577 40600 645697
rect 40000 645321 40600 645440
rect 677000 645245 677600 645311
rect 40000 645066 40600 645186
rect 677000 645106 677600 645172
rect 677000 644479 677600 644545
rect 677000 644309 677600 644375
rect 677000 644139 677600 644205
rect 40300 642252 40600 642322
rect 40300 641802 40600 641872
rect 677000 640328 677300 640398
rect 677000 639878 677300 639948
rect 40000 637995 40600 638061
rect 40000 637825 40600 637891
rect 40000 637655 40600 637721
rect 40000 637028 40600 637094
rect 677000 637014 677600 637134
rect 40000 636889 40600 636955
rect 677000 636760 677600 636879
rect 677000 636503 677600 636623
rect 677000 635927 677600 636047
rect 677000 635712 677600 635778
rect 677000 635511 677600 635577
rect 677000 635380 677600 635446
rect 40000 635058 40600 635178
rect 40000 633679 40600 633745
rect 40000 633509 40600 633575
rect 677000 633207 677600 633273
rect 677000 633058 677600 633124
rect 677000 632707 677600 632773
rect 677000 632258 677600 632324
rect 677000 631663 677600 631729
rect 40000 631169 40600 631243
rect 40000 629533 40600 629599
rect 40000 629363 40600 629429
rect 677000 628327 677600 628393
rect 677000 628063 677600 628129
rect 677000 627893 677600 627959
rect 40000 626825 40600 626891
rect 677000 626803 677600 626869
rect 40000 625387 40600 625453
rect 40000 625217 40600 625283
rect 40000 625047 40600 625113
rect 677000 624087 677600 624153
rect 677000 623917 677600 623983
rect 677000 623747 677600 623813
rect 40000 622331 40600 622397
rect 677000 622309 677600 622375
rect 40000 621241 40600 621307
rect 40000 621071 40600 621137
rect 40000 620807 40600 620873
rect 677000 619771 677600 619837
rect 677000 619601 677600 619667
rect 677000 617957 677600 618031
rect 40000 617471 40600 617537
rect 40000 616876 40600 616942
rect 40000 616427 40600 616493
rect 40000 616076 40600 616142
rect 40000 615927 40600 615993
rect 677000 615625 677600 615691
rect 677000 615455 677600 615521
rect 677000 614022 677600 614142
rect 40000 613754 40600 613820
rect 40000 613623 40600 613689
rect 40000 613422 40600 613488
rect 40000 613153 40600 613273
rect 40000 612577 40600 612697
rect 40000 612321 40600 612440
rect 677000 612245 677600 612311
rect 40000 612066 40600 612186
rect 677000 612106 677600 612172
rect 677000 611479 677600 611545
rect 677000 611309 677600 611375
rect 677000 611139 677600 611205
rect 40300 609252 40600 609322
rect 40300 608802 40600 608872
rect 677000 607328 677300 607398
rect 677000 606878 677300 606948
rect 40000 604995 40600 605061
rect 40000 604825 40600 604891
rect 40000 604655 40600 604721
rect 40000 604028 40600 604094
rect 677000 604014 677600 604134
rect 40000 603889 40600 603955
rect 677000 603760 677600 603879
rect 677000 603503 677600 603623
rect 677000 602927 677600 603047
rect 677000 602712 677600 602778
rect 677000 602511 677600 602577
rect 677000 602380 677600 602446
rect 40000 602058 40600 602178
rect 40000 600679 40600 600745
rect 40000 600509 40600 600575
rect 677000 600207 677600 600273
rect 677000 600058 677600 600124
rect 677000 599707 677600 599773
rect 677000 599258 677600 599324
rect 677000 598663 677600 598729
rect 40000 598169 40600 598243
rect 40000 596533 40600 596599
rect 40000 596363 40600 596429
rect 677000 595327 677600 595393
rect 677000 595063 677600 595129
rect 677000 594893 677600 594959
rect 40000 593825 40600 593891
rect 677000 593803 677600 593869
rect 40000 592387 40600 592453
rect 40000 592217 40600 592283
rect 40000 592047 40600 592113
rect 677000 591087 677600 591153
rect 677000 590917 677600 590983
rect 677000 590747 677600 590813
rect 40000 589331 40600 589397
rect 677000 589309 677600 589375
rect 40000 588241 40600 588307
rect 40000 588071 40600 588137
rect 40000 587807 40600 587873
rect 677000 586771 677600 586837
rect 677000 586601 677600 586667
rect 677000 584957 677600 585031
rect 40000 584471 40600 584537
rect 40000 583876 40600 583942
rect 40000 583427 40600 583493
rect 40000 583076 40600 583142
rect 40000 582927 40600 582993
rect 677000 582625 677600 582691
rect 677000 582455 677600 582521
rect 677000 581022 677600 581142
rect 40000 580754 40600 580820
rect 40000 580623 40600 580689
rect 40000 580422 40600 580488
rect 40000 580153 40600 580273
rect 40000 579577 40600 579697
rect 40000 579321 40600 579440
rect 677000 579245 677600 579311
rect 40000 579066 40600 579186
rect 677000 579106 677600 579172
rect 677000 578479 677600 578545
rect 677000 578309 677600 578375
rect 677000 578139 677600 578205
rect 40300 576252 40600 576322
rect 40300 575802 40600 575872
rect 677000 574328 677300 574398
rect 677000 573878 677300 573948
rect 40000 571995 40600 572061
rect 40000 571825 40600 571891
rect 40000 571655 40600 571721
rect 40000 571028 40600 571094
rect 677000 571014 677600 571134
rect 40000 570889 40600 570955
rect 677000 570760 677600 570879
rect 677000 570503 677600 570623
rect 677000 569927 677600 570047
rect 677000 569712 677600 569778
rect 677000 569511 677600 569577
rect 677000 569380 677600 569446
rect 40000 569058 40600 569178
rect 40000 567679 40600 567745
rect 40000 567509 40600 567575
rect 677000 567207 677600 567273
rect 677000 567058 677600 567124
rect 677000 566707 677600 566773
rect 677000 566258 677600 566324
rect 677000 565663 677600 565729
rect 40000 565169 40600 565243
rect 40000 563533 40600 563599
rect 40000 563363 40600 563429
rect 677000 562327 677600 562393
rect 677000 562063 677600 562129
rect 677000 561893 677600 561959
rect 40000 560825 40600 560891
rect 677000 560803 677600 560869
rect 40000 559387 40600 559453
rect 40000 559217 40600 559283
rect 40000 559047 40600 559113
rect 677000 558087 677600 558153
rect 677000 557917 677600 557983
rect 677000 557747 677600 557813
rect 40000 556331 40600 556397
rect 677000 556309 677600 556375
rect 40000 555241 40600 555307
rect 40000 555071 40600 555137
rect 40000 554807 40600 554873
rect 677000 553771 677600 553837
rect 677000 553601 677600 553667
rect 677000 551957 677600 552031
rect 40000 551471 40600 551537
rect 40000 550876 40600 550942
rect 40000 550427 40600 550493
rect 40000 550076 40600 550142
rect 40000 549927 40600 549993
rect 677000 549625 677600 549691
rect 677000 549455 677600 549521
rect 677000 548022 677600 548142
rect 40000 547754 40600 547820
rect 40000 547623 40600 547689
rect 40000 547422 40600 547488
rect 40000 547153 40600 547273
rect 40000 546577 40600 546697
rect 40000 546321 40600 546440
rect 677000 546245 677600 546311
rect 40000 546066 40600 546186
rect 677000 546106 677600 546172
rect 677000 545479 677600 545545
rect 677000 545309 677600 545375
rect 677000 545139 677600 545205
rect 677000 541328 677300 541398
rect 677000 540878 677300 540948
rect 39593 536078 40793 540858
rect 676807 533321 678007 538101
rect 39593 526099 40793 530879
rect 676807 523342 678007 528122
rect 27464 520530 28352 520570
rect 27464 517726 27504 520530
rect 28312 517726 28352 520530
rect 40000 518895 40600 519295
rect 27464 517686 28352 517726
rect 689246 517730 690136 517770
rect 677000 516161 677600 516561
rect 689246 514926 689286 517730
rect 690096 514926 690136 517730
rect 689246 514886 690136 514926
rect 40300 514476 40900 514536
rect 676700 513565 677300 513625
rect 40300 513495 40900 513555
rect 676700 513313 677300 513373
rect 40300 508897 40900 509025
rect 676700 508485 677300 508545
rect 40300 508141 40900 508201
rect 676700 508197 677300 508257
rect 40300 507943 40900 508003
rect 676700 507997 677300 508057
rect 40300 507743 40900 507803
rect 676700 507799 677300 507859
rect 40300 507455 40900 507515
rect 676700 506975 677300 507103
rect 40300 502627 40900 502687
rect 676700 502445 677300 502505
rect 40300 502375 40900 502435
rect 676700 501464 677300 501524
rect 39593 491551 40793 496340
rect 39593 489076 40793 491251
rect 39793 488776 40793 489076
rect 39593 486600 40793 488776
rect 676807 488700 678007 493502
rect 39593 481500 40793 486300
rect 676807 483748 677807 488410
rect 40300 478652 40600 478722
rect 676807 478660 678007 483449
rect 40300 478202 40600 478272
rect 40000 474395 40600 474461
rect 40000 474225 40600 474291
rect 40000 474055 40600 474121
rect 40000 473428 40600 473494
rect 677000 473414 677600 473534
rect 40000 473289 40600 473355
rect 677000 473160 677600 473279
rect 677000 472903 677600 473023
rect 677000 472327 677600 472447
rect 677000 472112 677600 472178
rect 677000 471911 677600 471977
rect 677000 471780 677600 471846
rect 40000 471458 40600 471578
rect 40000 470079 40600 470145
rect 40000 469909 40600 469975
rect 677000 469607 677600 469673
rect 677000 469458 677600 469524
rect 677000 469107 677600 469173
rect 677000 468658 677600 468724
rect 677000 468063 677600 468129
rect 40000 467569 40600 467643
rect 40000 465933 40600 465999
rect 40000 465763 40600 465829
rect 677000 464727 677600 464793
rect 677000 464463 677600 464529
rect 677000 464293 677600 464359
rect 40000 463225 40600 463291
rect 677000 463203 677600 463269
rect 40000 461787 40600 461853
rect 40000 461617 40600 461683
rect 40000 461447 40600 461513
rect 677000 460487 677600 460553
rect 677000 460317 677600 460383
rect 677000 460147 677600 460213
rect 40000 458731 40600 458797
rect 677000 458709 677600 458775
rect 40000 457641 40600 457707
rect 40000 457471 40600 457537
rect 40000 457207 40600 457273
rect 677000 456171 677600 456237
rect 677000 456001 677600 456067
rect 677000 454357 677600 454431
rect 40000 453871 40600 453937
rect 40000 453276 40600 453342
rect 40000 452827 40600 452893
rect 40000 452476 40600 452542
rect 40000 452327 40600 452393
rect 677000 452025 677600 452091
rect 677000 451855 677600 451921
rect 677000 450422 677600 450542
rect 40000 450154 40600 450220
rect 40000 450023 40600 450089
rect 40000 449822 40600 449888
rect 40000 449553 40600 449673
rect 40000 448977 40600 449097
rect 40000 448721 40600 448840
rect 677000 448645 677600 448711
rect 40000 448466 40600 448586
rect 677000 448506 677600 448572
rect 677000 447879 677600 447945
rect 677000 447709 677600 447775
rect 677000 447539 677600 447605
rect 40300 445652 40600 445722
rect 40300 445202 40600 445272
rect 677000 443728 677300 443798
rect 677000 443278 677300 443348
rect 40000 441395 40600 441461
rect 40000 441225 40600 441291
rect 40000 441055 40600 441121
rect 40000 440428 40600 440494
rect 677000 440414 677600 440534
rect 40000 440289 40600 440355
rect 677000 440160 677600 440279
rect 677000 439903 677600 440023
rect 677000 439327 677600 439447
rect 677000 439112 677600 439178
rect 677000 438911 677600 438977
rect 677000 438780 677600 438846
rect 40000 438458 40600 438578
rect 40000 437079 40600 437145
rect 40000 436909 40600 436975
rect 677000 436607 677600 436673
rect 677000 436458 677600 436524
rect 677000 436107 677600 436173
rect 677000 435658 677600 435724
rect 677000 435063 677600 435129
rect 40000 434569 40600 434643
rect 40000 432933 40600 432999
rect 40000 432763 40600 432829
rect 677000 431727 677600 431793
rect 677000 431463 677600 431529
rect 677000 431293 677600 431359
rect 40000 430225 40600 430291
rect 677000 430203 677600 430269
rect 40000 428787 40600 428853
rect 40000 428617 40600 428683
rect 40000 428447 40600 428513
rect 677000 427487 677600 427553
rect 677000 427317 677600 427383
rect 677000 427147 677600 427213
rect 40000 425731 40600 425797
rect 677000 425709 677600 425775
rect 40000 424641 40600 424707
rect 40000 424471 40600 424537
rect 40000 424207 40600 424273
rect 677000 423171 677600 423237
rect 677000 423001 677600 423067
rect 677000 421357 677600 421431
rect 40000 420871 40600 420937
rect 40000 420276 40600 420342
rect 40000 419827 40600 419893
rect 40000 419476 40600 419542
rect 40000 419327 40600 419393
rect 677000 419025 677600 419091
rect 677000 418855 677600 418921
rect 677000 417422 677600 417542
rect 40000 417154 40600 417220
rect 40000 417023 40600 417089
rect 40000 416822 40600 416888
rect 40000 416553 40600 416673
rect 40000 415977 40600 416097
rect 40000 415721 40600 415840
rect 677000 415645 677600 415711
rect 40000 415466 40600 415586
rect 677000 415506 677600 415572
rect 677000 414879 677600 414945
rect 677000 414709 677600 414775
rect 677000 414539 677600 414605
rect 40300 412652 40600 412722
rect 40300 412202 40600 412272
rect 677000 410728 677300 410798
rect 677000 410278 677300 410348
rect 40000 408395 40600 408461
rect 40000 408225 40600 408291
rect 40000 408055 40600 408121
rect 40000 407428 40600 407494
rect 677000 407414 677600 407534
rect 40000 407289 40600 407355
rect 677000 407160 677600 407279
rect 677000 406903 677600 407023
rect 677000 406327 677600 406447
rect 677000 406112 677600 406178
rect 677000 405911 677600 405977
rect 677000 405780 677600 405846
rect 40000 405458 40600 405578
rect 40000 404079 40600 404145
rect 40000 403909 40600 403975
rect 677000 403607 677600 403673
rect 677000 403458 677600 403524
rect 677000 403107 677600 403173
rect 677000 402658 677600 402724
rect 677000 402063 677600 402129
rect 40000 401569 40600 401643
rect 40000 399933 40600 399999
rect 40000 399763 40600 399829
rect 677000 398727 677600 398793
rect 677000 398463 677600 398529
rect 677000 398293 677600 398359
rect 40000 397225 40600 397291
rect 677000 397203 677600 397269
rect 40000 395787 40600 395853
rect 40000 395617 40600 395683
rect 40000 395447 40600 395513
rect 677000 394487 677600 394553
rect 677000 394317 677600 394383
rect 677000 394147 677600 394213
rect 40000 392731 40600 392797
rect 677000 392709 677600 392775
rect 40000 391641 40600 391707
rect 40000 391471 40600 391537
rect 40000 391207 40600 391273
rect 677000 390171 677600 390237
rect 677000 390001 677600 390067
rect 677000 388357 677600 388431
rect 40000 387871 40600 387937
rect 40000 387276 40600 387342
rect 40000 386827 40600 386893
rect 40000 386476 40600 386542
rect 40000 386327 40600 386393
rect 677000 386025 677600 386091
rect 677000 385855 677600 385921
rect 677000 384422 677600 384542
rect 40000 384154 40600 384220
rect 40000 384023 40600 384089
rect 40000 383822 40600 383888
rect 40000 383553 40600 383673
rect 40000 382977 40600 383097
rect 40000 382721 40600 382840
rect 677000 382645 677600 382711
rect 40000 382466 40600 382586
rect 677000 382506 677600 382572
rect 677000 381879 677600 381945
rect 677000 381709 677600 381775
rect 677000 381539 677600 381605
rect 40300 379652 40600 379722
rect 40300 379202 40600 379272
rect 677000 377728 677300 377798
rect 677000 377278 677300 377348
rect 40000 375395 40600 375461
rect 40000 375225 40600 375291
rect 40000 375055 40600 375121
rect 40000 374428 40600 374494
rect 677000 374414 677600 374534
rect 40000 374289 40600 374355
rect 677000 374160 677600 374279
rect 677000 373903 677600 374023
rect 677000 373327 677600 373447
rect 677000 373112 677600 373178
rect 677000 372911 677600 372977
rect 677000 372780 677600 372846
rect 40000 372458 40600 372578
rect 40000 371079 40600 371145
rect 40000 370909 40600 370975
rect 677000 370607 677600 370673
rect 677000 370458 677600 370524
rect 677000 370107 677600 370173
rect 677000 369658 677600 369724
rect 677000 369063 677600 369129
rect 40000 368569 40600 368643
rect 40000 366933 40600 366999
rect 40000 366763 40600 366829
rect 677000 365727 677600 365793
rect 677000 365463 677600 365529
rect 677000 365293 677600 365359
rect 40000 364225 40600 364291
rect 677000 364203 677600 364269
rect 40000 362787 40600 362853
rect 40000 362617 40600 362683
rect 40000 362447 40600 362513
rect 677000 361487 677600 361553
rect 677000 361317 677600 361383
rect 677000 361147 677600 361213
rect 40000 359731 40600 359797
rect 677000 359709 677600 359775
rect 40000 358641 40600 358707
rect 40000 358471 40600 358537
rect 40000 358207 40600 358273
rect 677000 357171 677600 357237
rect 677000 357001 677600 357067
rect 677000 355357 677600 355431
rect 40000 354871 40600 354937
rect 40000 354276 40600 354342
rect 40000 353827 40600 353893
rect 40000 353476 40600 353542
rect 40000 353327 40600 353393
rect 677000 353025 677600 353091
rect 677000 352855 677600 352921
rect 677000 351422 677600 351542
rect 40000 351154 40600 351220
rect 40000 351023 40600 351089
rect 40000 350822 40600 350888
rect 40000 350553 40600 350673
rect 40000 349977 40600 350097
rect 40000 349721 40600 349840
rect 677000 349645 677600 349711
rect 40000 349466 40600 349586
rect 677000 349506 677600 349572
rect 677000 348879 677600 348945
rect 677000 348709 677600 348775
rect 677000 348539 677600 348605
rect 677000 344728 677300 344798
rect 677000 344278 677300 344348
rect 39593 339478 40793 344258
rect 676807 336721 678007 341501
rect 39593 329499 40793 334279
rect 676807 326742 678007 331522
rect 39593 316478 40793 321258
rect 676807 312721 678007 317501
rect 39593 306499 40793 311279
rect 676807 302742 678007 307522
rect 39593 296478 40793 301258
rect 676807 292721 678007 297501
rect 39593 286499 40793 291279
rect 40542 283652 40842 283722
rect 40542 283202 40842 283272
rect 676807 282742 678007 287522
rect 40542 282002 40842 282072
rect 40542 281704 40842 281774
rect 40538 281424 40838 281494
rect 40542 281112 40842 281182
rect 40542 280838 40842 280908
rect 40542 280490 40842 280618
rect 40542 279058 40842 279188
rect 40542 278528 40842 278598
rect 40542 277964 40842 278178
rect 40542 277332 40842 277402
rect 676758 277396 677058 277520
rect 676758 276868 677058 276938
rect 676758 276458 677058 276528
rect 676758 276114 677058 276184
rect 676758 275252 677058 275322
rect 40542 275120 40842 275190
rect 40542 274572 40842 274642
rect 676758 274532 677058 274602
rect 40542 273992 40842 274062
rect 676758 273332 677058 273402
rect 40542 272826 40842 272896
rect 676758 272560 677058 272630
rect 40542 272370 40842 272440
rect 676758 272076 677058 272146
rect 40542 271916 40842 271986
rect 676758 271632 677058 271702
rect 40542 271298 40842 271368
rect 676758 271014 677058 271084
rect 40542 270854 40842 270924
rect 676758 270560 677058 270630
rect 40542 270370 40842 270440
rect 676758 270104 677058 270174
rect 40542 269598 40842 269668
rect 676758 268938 677058 269008
rect 40542 268398 40842 268468
rect 676758 268358 677058 268428
rect 676758 267810 677058 267880
rect 40542 267678 40842 267748
rect 40542 266816 40842 266886
rect 40542 266472 40842 266542
rect 40542 266062 40842 266132
rect 40542 265480 40842 265604
rect 676758 265598 677058 265668
rect 676758 264822 677058 265036
rect 676758 264402 677058 264472
rect 676758 263812 677058 263942
rect 40542 262652 40842 262722
rect 676758 262382 677058 262510
rect 40542 262202 40842 262272
rect 676758 262092 677058 262162
rect 676758 261818 677058 261888
rect 676762 261506 677062 261576
rect 676758 261226 677058 261296
rect 40542 261002 40842 261072
rect 676758 260928 677058 260998
rect 40542 260704 40842 260774
rect 40538 260424 40838 260494
rect 40542 260112 40842 260182
rect 40542 259838 40842 259908
rect 676758 259728 677058 259798
rect 40542 259490 40842 259618
rect 676758 259278 677058 259348
rect 40542 258058 40842 258188
rect 40542 257528 40842 257598
rect 40542 256964 40842 257178
rect 40542 256332 40842 256402
rect 676758 256396 677058 256520
rect 676758 255868 677058 255938
rect 676758 255458 677058 255528
rect 676758 255114 677058 255184
rect 676758 254252 677058 254322
rect 40542 254120 40842 254190
rect 40542 253572 40842 253642
rect 676758 253532 677058 253602
rect 40542 252992 40842 253062
rect 676758 252332 677058 252402
rect 40542 251826 40842 251896
rect 676758 251560 677058 251630
rect 40542 251370 40842 251440
rect 676758 251076 677058 251146
rect 40542 250916 40842 250986
rect 676758 250632 677058 250702
rect 40542 250298 40842 250368
rect 676758 250014 677058 250084
rect 40542 249854 40842 249924
rect 676758 249560 677058 249630
rect 40542 249370 40842 249440
rect 676758 249104 677058 249174
rect 40542 248598 40842 248668
rect 676758 247938 677058 248008
rect 40542 247398 40842 247468
rect 676758 247358 677058 247428
rect 676758 246810 677058 246880
rect 40542 246678 40842 246748
rect 40542 245816 40842 245886
rect 40542 245472 40842 245542
rect 40542 245062 40842 245132
rect 40542 244480 40842 244604
rect 676758 244598 677058 244668
rect 676758 243822 677058 244036
rect 676758 243402 677058 243472
rect 676758 242812 677058 242942
rect 40542 241652 40842 241722
rect 676758 241382 677058 241510
rect 40542 241202 40842 241272
rect 676758 241092 677058 241162
rect 676758 240818 677058 240888
rect 676762 240506 677062 240576
rect 676758 240226 677058 240296
rect 40542 240002 40842 240072
rect 676758 239928 677058 239998
rect 40542 239704 40842 239774
rect 40538 239424 40838 239494
rect 40542 239112 40842 239182
rect 40542 238838 40842 238908
rect 676758 238728 677058 238798
rect 40542 238490 40842 238618
rect 676758 238278 677058 238348
rect 40542 237058 40842 237188
rect 40542 236528 40842 236598
rect 40542 235964 40842 236178
rect 40542 235332 40842 235402
rect 676758 235396 677058 235520
rect 676758 234868 677058 234938
rect 676758 234458 677058 234528
rect 676758 234114 677058 234184
rect 676758 233252 677058 233322
rect 40542 233120 40842 233190
rect 40542 232572 40842 232642
rect 676758 232532 677058 232602
rect 40542 231992 40842 232062
rect 676758 231332 677058 231402
rect 40542 230826 40842 230896
rect 676758 230560 677058 230630
rect 40542 230370 40842 230440
rect 676758 230076 677058 230146
rect 40542 229916 40842 229986
rect 676758 229632 677058 229702
rect 40542 229298 40842 229368
rect 676758 229014 677058 229084
rect 40542 228854 40842 228924
rect 676758 228560 677058 228630
rect 40542 228370 40842 228440
rect 676758 228104 677058 228174
rect 40542 227598 40842 227668
rect 676758 226938 677058 227008
rect 40542 226398 40842 226468
rect 676758 226358 677058 226428
rect 676758 225810 677058 225880
rect 40542 225678 40842 225748
rect 40542 224816 40842 224886
rect 40542 224472 40842 224542
rect 40542 224062 40842 224132
rect 40542 223480 40842 223604
rect 676758 223598 677058 223668
rect 676758 222822 677058 223036
rect 676758 222402 677058 222472
rect 676758 221812 677058 221942
rect 40542 220652 40842 220722
rect 676758 220382 677058 220510
rect 40542 220202 40842 220272
rect 676758 220092 677058 220162
rect 676758 219818 677058 219888
rect 676762 219506 677062 219576
rect 676758 219226 677058 219296
rect 40542 219002 40842 219072
rect 676758 218928 677058 218998
rect 40542 218704 40842 218774
rect 40538 218424 40838 218494
rect 40542 218112 40842 218182
rect 40542 217838 40842 217908
rect 676758 217728 677058 217798
rect 40542 217490 40842 217618
rect 676758 217278 677058 217348
rect 40542 216058 40842 216188
rect 40542 215528 40842 215598
rect 40542 214964 40842 215178
rect 40542 214332 40842 214402
rect 676758 214396 677058 214520
rect 676758 213868 677058 213938
rect 676758 213458 677058 213528
rect 676758 213114 677058 213184
rect 676758 212252 677058 212322
rect 40542 212120 40842 212190
rect 40542 211572 40842 211642
rect 676758 211532 677058 211602
rect 40542 210992 40842 211062
rect 676758 210332 677058 210402
rect 40542 209826 40842 209896
rect 676758 209560 677058 209630
rect 40542 209370 40842 209440
rect 676758 209076 677058 209146
rect 40542 208916 40842 208986
rect 676758 208632 677058 208702
rect 40542 208298 40842 208368
rect 676758 208014 677058 208084
rect 40542 207854 40842 207924
rect 676758 207560 677058 207630
rect 40542 207370 40842 207440
rect 676758 207104 677058 207174
rect 40542 206598 40842 206668
rect 676758 205938 677058 206008
rect 40542 205398 40842 205468
rect 676758 205358 677058 205428
rect 676758 204810 677058 204880
rect 40542 204678 40842 204748
rect 40542 203816 40842 203886
rect 40542 203472 40842 203542
rect 40542 203062 40842 203132
rect 40542 202480 40842 202604
rect 676758 202598 677058 202668
rect 676758 201822 677058 202036
rect 676758 201402 677058 201472
rect 676758 200812 677058 200942
rect 676758 199382 677058 199510
rect 676758 199092 677058 199162
rect 676758 198818 677058 198888
rect 676762 198506 677062 198576
rect 676758 198226 677058 198296
rect 676758 197928 677058 197998
rect 39593 192478 40793 197258
rect 676758 196728 677058 196798
rect 676758 196278 677058 196348
rect 676807 188721 678007 193501
rect 39593 182499 40793 187279
rect 676807 178742 678007 183522
rect 39593 169551 40793 174340
rect 39793 164590 40793 169252
rect 676807 168700 678007 173500
rect 676807 166224 678007 168400
rect 676807 165924 677807 166224
rect 39593 159498 40793 164300
rect 676807 163749 678007 165924
rect 676807 158660 678007 163449
rect 40542 156652 40842 156722
rect 40542 156202 40842 156272
rect 40542 155002 40842 155072
rect 40542 154704 40842 154774
rect 40538 154424 40838 154494
rect 40542 154112 40842 154182
rect 40542 153838 40842 153908
rect 40542 153490 40842 153618
rect 676758 153396 677058 153520
rect 676758 152868 677058 152938
rect 676758 152458 677058 152528
rect 40542 152058 40842 152188
rect 676758 152114 677058 152184
rect 40542 151528 40842 151598
rect 676758 151252 677058 151322
rect 40542 150964 40842 151178
rect 676758 150532 677058 150602
rect 40542 150332 40842 150402
rect 676758 149332 677058 149402
rect 676758 148560 677058 148630
rect 40542 148120 40842 148190
rect 676758 148076 677058 148146
rect 40542 147572 40842 147642
rect 676758 147632 677058 147702
rect 40542 146992 40842 147062
rect 676758 147014 677058 147084
rect 676758 146560 677058 146630
rect 676758 146104 677058 146174
rect 40542 145826 40842 145896
rect 40542 145370 40842 145440
rect 40542 144916 40842 144986
rect 676758 144938 677058 145008
rect 40542 144298 40842 144368
rect 676758 144358 677058 144428
rect 40542 143854 40842 143924
rect 676758 143810 677058 143880
rect 40542 143370 40842 143440
rect 40542 142598 40842 142668
rect 676758 141598 677058 141668
rect 40542 141398 40842 141468
rect 676758 140822 677058 141036
rect 40542 140678 40842 140748
rect 676758 140402 677058 140472
rect 40542 139816 40842 139886
rect 676758 139812 677058 139942
rect 40542 139472 40842 139542
rect 40542 139062 40842 139132
rect 40542 138480 40842 138604
rect 676758 138382 677058 138510
rect 676758 138092 677058 138162
rect 676758 137818 677058 137888
rect 676762 137506 677062 137576
rect 676758 137226 677058 137296
rect 676758 136928 677058 136998
rect 676758 135728 677058 135798
rect 40542 135652 40842 135722
rect 676758 135278 677058 135348
rect 40542 135202 40842 135272
rect 40542 134002 40842 134072
rect 40542 133704 40842 133774
rect 40538 133424 40838 133494
rect 40542 133112 40842 133182
rect 40542 132838 40842 132908
rect 40542 132490 40842 132618
rect 676758 132396 677058 132520
rect 676758 131868 677058 131938
rect 676758 131458 677058 131528
rect 40542 131058 40842 131188
rect 676758 131114 677058 131184
rect 40542 130528 40842 130598
rect 676758 130252 677058 130322
rect 40542 129964 40842 130178
rect 676758 129532 677058 129602
rect 40542 129332 40842 129402
rect 676758 128332 677058 128402
rect 676758 127560 677058 127630
rect 40542 127120 40842 127190
rect 676758 127076 677058 127146
rect 40542 126572 40842 126642
rect 676758 126632 677058 126702
rect 40542 125992 40842 126062
rect 676758 126014 677058 126084
rect 676758 125560 677058 125630
rect 676758 125104 677058 125174
rect 40542 124826 40842 124896
rect 40542 124370 40842 124440
rect 40542 123916 40842 123986
rect 676758 123938 677058 124008
rect 40542 123298 40842 123368
rect 676758 123358 677058 123428
rect 40542 122854 40842 122924
rect 676758 122810 677058 122880
rect 40542 122370 40842 122440
rect 40542 121598 40842 121668
rect 676758 120598 677058 120668
rect 40542 120398 40842 120468
rect 676758 119822 677058 120036
rect 40542 119678 40842 119748
rect 676758 119402 677058 119472
rect 40542 118816 40842 118886
rect 676758 118812 677058 118942
rect 40542 118472 40842 118542
rect 40542 118062 40842 118132
rect 40542 117480 40842 117604
rect 676758 117382 677058 117510
rect 676758 117092 677058 117162
rect 676758 116818 677058 116888
rect 676762 116506 677062 116576
rect 676758 116226 677058 116296
rect 676758 115928 677058 115998
rect 676758 114728 677058 114798
rect 40542 114652 40842 114722
rect 676758 114278 677058 114348
rect 40542 114202 40842 114272
rect 40542 113002 40842 113072
rect 40542 112704 40842 112774
rect 40538 112424 40838 112494
rect 40542 112112 40842 112182
rect 40542 111838 40842 111908
rect 40542 111490 40842 111618
rect 676758 111396 677058 111520
rect 676758 110868 677058 110938
rect 676758 110458 677058 110528
rect 40542 110058 40842 110188
rect 676758 110114 677058 110184
rect 40542 109528 40842 109598
rect 676758 109252 677058 109322
rect 40542 108964 40842 109178
rect 676758 108532 677058 108602
rect 40542 108332 40842 108402
rect 676758 107332 677058 107402
rect 676758 106560 677058 106630
rect 40542 106120 40842 106190
rect 676758 106076 677058 106146
rect 40542 105572 40842 105642
rect 676758 105632 677058 105702
rect 40542 104992 40842 105062
rect 676758 105014 677058 105084
rect 676758 104560 677058 104630
rect 676758 104104 677058 104174
rect 40542 103826 40842 103896
rect 40542 103370 40842 103440
rect 40542 102916 40842 102986
rect 676758 102938 677058 103008
rect 40542 102298 40842 102368
rect 676758 102358 677058 102428
rect 40542 101854 40842 101924
rect 676758 101810 677058 101880
rect 40542 101370 40842 101440
rect 40542 100598 40842 100668
rect 676758 99598 677058 99668
rect 40542 99398 40842 99468
rect 676758 98822 677058 99036
rect 40542 98678 40842 98748
rect 676758 98402 677058 98472
rect 40542 97816 40842 97886
rect 676758 97812 677058 97942
rect 40542 97472 40842 97542
rect 40542 97062 40842 97132
rect 40542 96480 40842 96604
rect 676758 96382 677058 96510
rect 676758 96092 677058 96162
rect 676758 95818 677058 95888
rect 676762 95506 677062 95576
rect 676758 95226 677058 95296
rect 676758 94928 677058 94998
rect 676758 93728 677058 93798
rect 40542 93652 40842 93722
rect 676758 93278 677058 93348
rect 40542 93202 40842 93272
rect 40542 92002 40842 92072
rect 40542 91704 40842 91774
rect 40538 91424 40838 91494
rect 40542 91112 40842 91182
rect 40542 90838 40842 90908
rect 40542 90490 40842 90618
rect 676758 90396 677058 90520
rect 676758 89868 677058 89938
rect 676758 89458 677058 89528
rect 40542 89058 40842 89188
rect 676758 89114 677058 89184
rect 40542 88528 40842 88598
rect 676758 88252 677058 88322
rect 40542 87964 40842 88178
rect 676758 87532 677058 87602
rect 40542 87332 40842 87402
rect 676758 86332 677058 86402
rect 676758 85560 677058 85630
rect 40542 85120 40842 85190
rect 676758 85076 677058 85146
rect 40542 84572 40842 84642
rect 676758 84632 677058 84702
rect 40542 83992 40842 84062
rect 676758 84014 677058 84084
rect 676758 83560 677058 83630
rect 676758 83104 677058 83174
rect 40542 82826 40842 82896
rect 40542 82370 40842 82440
rect 40542 81916 40842 81986
rect 676758 81938 677058 82008
rect 40542 81298 40842 81368
rect 676758 81358 677058 81428
rect 40542 80854 40842 80924
rect 676758 80810 677058 80880
rect 40542 80370 40842 80440
rect 40542 79598 40842 79668
rect 676758 78598 677058 78668
rect 40542 78398 40842 78468
rect 676758 77822 677058 78036
rect 40542 77678 40842 77748
rect 676758 77402 677058 77472
rect 40542 76816 40842 76886
rect 676758 76812 677058 76942
rect 40542 76472 40842 76542
rect 40542 76062 40842 76132
rect 40542 75480 40842 75604
rect 676758 75382 677058 75510
rect 676758 75092 677058 75162
rect 676758 74818 677058 74888
rect 676762 74506 677062 74576
rect 676758 74226 677058 74296
rect 676758 73928 677058 73998
rect 676758 72728 677058 72798
rect 676758 72278 677058 72348
rect 39593 65478 40793 70258
rect 676807 64721 678007 69501
rect 39593 55499 40793 60279
rect 676807 54742 678007 59522
rect 676700 48232 677300 48292
rect 40300 47954 40900 48014
rect 676700 47896 677300 47956
rect 676700 47644 677300 47704
rect 676700 47392 677300 47452
rect 676700 47140 677300 47200
rect 40300 47074 40900 47134
rect 676700 46888 677300 46948
rect 40300 43452 40900 43512
rect 676700 43266 677300 43326
rect 40300 43200 40900 43260
rect 40300 42948 40900 43008
rect 40300 42696 40900 42756
rect 40300 42444 40900 42504
rect 676700 42386 677300 42446
rect 40300 42108 40900 42168
rect 47060 39593 51849 40793
rect 57100 39593 61902 40793
rect 206142 39593 210922 40793
rect 216121 39593 220901 40793
rect 228060 39593 232849 40793
rect 238100 39593 242900 40793
rect 255438 40388 257234 40400
rect 255438 40012 255450 40388
rect 257222 40012 257234 40388
rect 255438 39600 257234 40012
rect 277438 40388 279234 40400
rect 277438 40012 277450 40388
rect 279222 40012 279234 40388
rect 277438 39600 279234 40012
rect 299438 40388 301234 40400
rect 299438 40012 299450 40388
rect 301222 40012 301234 40388
rect 299438 39600 301234 40012
rect 321438 40388 323234 40400
rect 321438 40012 321450 40388
rect 323222 40012 323234 40388
rect 321438 39600 323234 40012
rect 338142 39593 342922 40793
rect 348121 39593 352901 40793
rect 364060 39593 368849 40793
rect 374100 39593 378902 40793
rect 478142 39593 482922 40793
rect 488121 39593 492901 40793
rect 500142 39593 504922 40793
rect 510121 39593 514901 40793
rect 526142 39593 530922 40793
rect 536121 39593 540901 40793
rect 552060 39593 556849 40793
rect 562100 39593 566900 40793
<< via3 >>
rect 27504 517726 28312 520530
rect 689286 514926 690096 517730
<< metal5 >>
rect 48300 1020680 56300 1028680
rect 72300 1020757 80300 1028757
rect 96300 1020757 104300 1028757
rect 120300 1020757 128300 1028757
rect 144300 1020757 152300 1028757
rect 167300 1020680 175300 1028680
rect 190300 1020680 198300 1028680
rect 214300 1020757 222300 1028757
rect 238300 1020757 246300 1028757
rect 262300 1020757 270300 1028757
rect 286300 1020757 294300 1028757
rect 309300 1020680 317300 1028680
rect 332300 1020680 340300 1028680
rect 355300 1020680 363300 1028680
rect 378300 1020680 386300 1028680
rect 401300 1020680 409300 1028680
rect 425300 1020757 433300 1028757
rect 449300 1020757 457300 1028757
rect 473300 1020757 481300 1028757
rect 497300 1020757 505300 1028757
rect 520300 1020680 528300 1028680
rect 543300 1020680 551300 1028680
rect 567300 1020757 575300 1028757
rect 591300 1020757 599300 1028757
rect 615300 1020757 623300 1028757
rect 639300 1020757 647300 1028757
rect 662300 1020680 670300 1028680
rect 8920 975500 16920 983500
rect 700680 974700 708680 982700
rect 8920 952500 16920 960500
rect 700680 950700 708680 958700
rect 8843 932500 16843 940500
rect 700757 929700 708757 937700
rect 8843 911500 16843 919500
rect 700757 908700 708757 916700
rect 8843 890500 16843 898500
rect 700757 887700 708757 895700
rect 8843 869500 16843 877500
rect 700757 866700 708757 874700
rect 8920 848500 16920 856500
rect 700680 846700 708680 854700
rect 8843 828500 16843 836500
rect 700757 825700 708757 833700
rect 8843 807500 16843 815500
rect 700757 804700 708757 812700
rect 8843 786500 16843 794500
rect 700757 783700 708757 791700
rect 8843 765500 16843 773500
rect 700757 762700 708757 770700
rect 8920 744500 16920 752500
rect 700680 742700 708680 750700
rect 8920 724500 16920 732500
rect 700680 722700 708680 730700
rect 8920 701500 16920 709500
rect 700680 698700 708680 706700
rect 8920 681500 16920 689500
rect 700680 678700 708680 686700
rect 8504 651866 16504 659866
rect 701096 655334 709096 663334
rect 8504 618866 16504 626866
rect 701096 622334 709096 630334
rect 8504 585866 16504 593866
rect 701096 589334 709096 597334
rect 8504 552866 16504 560866
rect 701096 556334 709096 564334
rect 8920 529500 16920 537500
rect 700680 526700 708680 534700
rect 8920 484900 16920 492900
rect 700680 482100 708680 490100
rect 8504 455266 16504 463266
rect 701096 458734 709096 466734
rect 8504 422266 16504 430266
rect 701096 425734 709096 433734
rect 8504 389266 16504 397266
rect 701096 392734 709096 400734
rect 8504 356266 16504 364266
rect 701096 359734 709096 367734
rect 8920 332900 16920 340900
rect 700680 330100 708680 338100
rect 8920 309900 16920 317900
rect 700680 306100 708680 314100
rect 8920 289900 16920 297900
rect 700680 286100 708680 294100
rect 8843 269900 16843 277900
rect 700757 265100 708757 273100
rect 8843 248900 16843 256900
rect 700757 244100 708757 252100
rect 8843 227900 16843 235900
rect 700757 223100 708757 231100
rect 8843 206900 16843 214900
rect 700757 202100 708757 210100
rect 8920 185900 16920 193900
rect 700680 182100 708680 190100
rect 8920 162900 16920 170900
rect 700680 162100 708680 170100
rect 8843 142900 16843 150900
rect 700757 141100 708757 149100
rect 8843 121900 16843 129900
rect 700757 120100 708757 128100
rect 8843 100900 16843 108900
rect 700757 99100 708757 107100
rect 8843 79900 16843 87900
rect 700757 78100 708757 86100
rect 8920 58900 16920 66900
rect 700680 58100 708680 66100
rect 50500 8920 58500 16920
rect 72500 8843 80500 16843
rect 95500 8920 103500 16920
rect 117500 8843 125500 16843
rect 140500 8843 148500 16843
rect 163500 8843 171500 16843
rect 186500 8843 194500 16843
rect 209500 8920 217500 16920
rect 231500 8920 239500 16920
rect 253500 8920 261500 16920
rect 275500 8920 283500 16920
rect 297500 8920 305500 16920
rect 319500 8920 327500 16920
rect 341500 8920 349500 16920
rect 367500 8920 375500 16920
rect 389500 8843 397500 16843
rect 412500 8843 420500 16843
rect 435500 8843 443500 16843
rect 458500 8843 466500 16843
rect 481500 8920 489500 16920
rect 503500 8920 511500 16920
rect 529500 8920 537500 16920
rect 555500 8920 563500 16920
rect 615697 14068 623697 22068
rect 638302 14068 646302 22068
use sky130_fd_io__top_analog_pad  analog_0_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 1 0 351800 0 1 998000
box -80 0 15080 39600
use sky130_fd_io__top_analog_pad  analog_1_pad
timestamp 1726580063
transform 1 0 328800 0 1 998000
box -80 0 15080 39600
use caravel_logo  caravel_logo_0
timestamp 1638586901
transform 1 0 6820 0 1 1007840
box -2520 0 15000 15560
use caravel_motto  caravel_motto_0
timestamp 1637698310
transform 1 0 -351120 0 1 1002542
box 373080 14838 395618 19242
use copyright_block_frigate  copyright_block_frigate_0
timestamp 1706137558
transform 1 0 671202 0 1 16828
box -262 -10348 30014 2764
use sky130_ef_io__corner_pad  corner_ne $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 1 0 677600 0 1 996800
box 0 0 40000 40800
use sky130_ef_io__corner_pad  corner_nw
timestamp 1726580063
transform 0 -1 40800 1 0 997600
box 0 0 40000 40800
use sky130_ef_io__corner_pad  corner_se
timestamp 1726580063
transform 0 1 676800 -1 0 40000
box 0 0 40000 40800
use sky130_ef_io__corner_pad  corner_sw
timestamp 1726580063
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use chip_io_gpio_connects_horiz  gpio0_0_connects
timestamp 1706150479
transform 1 0 676758 0 1 73830
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio0_0_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 0 1 678007 -1 0 90600
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio0_1_connects
timestamp 1706150479
transform 1 0 676758 0 1 94830
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio0_1_pad
timestamp 1726580063
transform 0 1 678007 -1 0 111600
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio0_2_connects
timestamp 1706150479
transform 1 0 676758 0 1 115830
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio0_2_pad
timestamp 1726580063
transform 0 1 678007 -1 0 132600
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio0_3_connects
timestamp 1706150479
transform 1 0 676758 0 1 136830
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio0_3_pad
timestamp 1726580063
transform 0 1 678007 -1 0 153600
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio0_4_connects
timestamp 1706150479
transform 1 0 676758 0 1 197830
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio0_4_pad
timestamp 1726580063
transform 0 1 678007 -1 0 214600
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio0_5_connects
timestamp 1706150479
transform 1 0 676758 0 1 218830
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio0_5_pad
timestamp 1726580063
transform 0 1 678007 -1 0 235600
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio0_6_connects
timestamp 1706150479
transform 1 0 676758 0 1 239830
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio0_6_pad
timestamp 1726580063
transform 0 1 678007 -1 0 256600
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio0_7_connects
timestamp 1706150479
transform 1 0 676758 0 1 260830
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio0_7_pad
timestamp 1726580063
transform 0 1 678007 -1 0 277600
box -143 -407 16134 39593
use chip_io_ovt_connects_horiz  gpio1_0_connects
timestamp 1706150479
transform 1 0 676760 0 1 345830
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio1_0_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 0 1 677600 -1 0 374600
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio1_1_connects
timestamp 1706150479
transform 1 0 676760 0 1 378830
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio1_1_pad
timestamp 1726580063
transform 0 1 677600 -1 0 407600
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio1_2_connects
timestamp 1706150479
transform 1 0 676760 0 1 411830
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio1_2_pad
timestamp 1726580063
transform 0 1 677600 -1 0 440600
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio1_3_connects
timestamp 1706150479
transform 1 0 676760 0 1 444830
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio1_3_pad
timestamp 1726580063
transform 0 1 677600 -1 0 473600
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio1_4_connects
timestamp 1706150479
transform 1 0 676760 0 1 542430
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio1_4_pad
timestamp 1726580063
transform 0 1 677600 -1 0 571200
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio1_5_connects
timestamp 1706150479
transform 1 0 676760 0 1 575430
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio1_5_pad
timestamp 1726580063
transform 0 1 677600 -1 0 604200
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio1_6_connects
timestamp 1706150479
transform 1 0 676760 0 1 608430
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio1_6_pad
timestamp 1726580063
transform 0 1 677600 -1 0 637200
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio1_7_connects
timestamp 1706150479
transform 1 0 676760 0 1 641430
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio1_7_pad
timestamp 1726580063
transform 0 1 677600 -1 0 670200
box -80 -147 28211 40151
use chip_io_gpio_connects_horiz  gpio2_0_connects
timestamp 1706150479
transform 1 0 676758 0 1 758430
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio2_0_pad
timestamp 1726580063
transform 0 1 678007 -1 0 775200
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio2_1_connects
timestamp 1706150479
transform 1 0 676758 0 1 779430
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio2_1_pad
timestamp 1726580063
transform 0 1 678007 -1 0 796200
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio2_2_connects
timestamp 1706150479
transform 1 0 676758 0 1 800430
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio2_2_pad
timestamp 1726580063
transform 0 1 678007 -1 0 817200
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio2_3_connects
timestamp 1706150479
transform 1 0 676758 0 1 821430
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio2_3_pad
timestamp 1726580063
transform 0 1 678007 -1 0 838200
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio2_4_connects
timestamp 1706150479
transform 1 0 676758 0 1 862430
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio2_4_pad
timestamp 1726580063
transform 0 1 678007 -1 0 879200
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio2_5_connects
timestamp 1706150479
transform 1 0 676758 0 1 883430
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio2_5_pad
timestamp 1726580063
transform 0 1 678007 -1 0 900200
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio2_6_connects
timestamp 1706150479
transform 1 0 676758 0 1 904430
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio2_6_pad
timestamp 1726580063
transform 0 1 678007 -1 0 921200
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio2_7_connects
timestamp 1706150479
transform 1 0 676758 0 1 925430
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio2_7_pad
timestamp 1726580063
transform 0 1 678007 -1 0 942200
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio3_0_connects
timestamp 1726510233
transform 0 -1 651456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio3_0_pad
timestamp 1726580063
transform 1 0 634800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio3_1_connects
timestamp 1726510233
transform 0 -1 627456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio3_1_pad
timestamp 1726580063
transform 1 0 610800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio3_2_connects
timestamp 1726510233
transform 0 -1 603456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio3_2_pad
timestamp 1726580063
transform 1 0 586800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio3_3_connects
timestamp 1726510233
transform 0 -1 579456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio3_3_pad
timestamp 1726580063
transform 1 0 562800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio3_4_connects
timestamp 1726510233
transform 0 -1 509456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio3_4_pad
timestamp 1726580063
transform 1 0 492800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio3_5_connects
timestamp 1726510233
transform 0 -1 485456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio3_5_pad
timestamp 1726580063
transform 1 0 468800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio3_6_connects
timestamp 1726510233
transform 0 -1 461456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio3_6_pad
timestamp 1726580063
transform 1 0 444800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio3_7_connects
timestamp 1726510233
transform 0 -1 437456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio3_7_pad
timestamp 1726580063
transform 1 0 420800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio4_0_connects
timestamp 1726510233
transform 0 -1 298456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio4_0_pad
timestamp 1726580063
transform 1 0 281800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio4_1_connects
timestamp 1726510233
transform 0 -1 274456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio4_1_pad
timestamp 1726580063
transform 1 0 257800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio4_2_connects
timestamp 1726510233
transform 0 -1 250456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio4_2_pad
timestamp 1726580063
transform 1 0 233800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio4_3_connects
timestamp 1726510233
transform 0 -1 226456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio4_3_pad
timestamp 1726580063
transform 1 0 209800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio4_4_connects
timestamp 1726510233
transform 0 -1 156456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio4_4_pad
timestamp 1726580063
transform 1 0 139800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio4_5_connects
timestamp 1726510233
transform 0 -1 132456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio4_5_pad
timestamp 1726580063
transform 1 0 115800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio4_6_connects
timestamp 1726510233
transform 0 -1 108456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio4_6_pad
timestamp 1726580063
transform 1 0 91800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio4_7_connects
timestamp 1726510233
transform 0 -1 84456 1 0 996690
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio4_7_pad
timestamp 1726580063
transform 1 0 67800 0 1 998007
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio5_0_connects
timestamp 1706150479
transform -1 0 40842 0 -1 944770
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio5_0_pad
timestamp 1726580063
transform 0 -1 39593 1 0 928000
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio5_1_connects
timestamp 1706150479
transform -1 0 40842 0 -1 923770
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio5_1_pad
timestamp 1726580063
transform 0 -1 39593 1 0 907000
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio5_2_connects
timestamp 1706150479
transform -1 0 40842 0 -1 902770
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio5_2_pad
timestamp 1726580063
transform 0 -1 39593 1 0 886000
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio5_3_connects
timestamp 1706150479
transform -1 0 40842 0 -1 881770
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio5_3_pad
timestamp 1726580063
transform 0 -1 39593 1 0 865000
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio5_4_connects
timestamp 1706150479
transform -1 0 40842 0 -1 840770
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio5_4_pad
timestamp 1726580063
transform 0 -1 39593 1 0 824000
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio5_5_connects
timestamp 1706150479
transform -1 0 40842 0 -1 819770
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio5_5_pad
timestamp 1726580063
transform 0 -1 39593 1 0 803000
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio5_6_connects
timestamp 1706150479
transform -1 0 40842 0 -1 798770
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio5_6_pad
timestamp 1726580063
transform 0 -1 39593 1 0 782000
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio5_7_connects
timestamp 1706150479
transform -1 0 40842 0 -1 777770
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio5_7_pad
timestamp 1726580063
transform 0 -1 39593 1 0 761000
box -143 -407 16134 39593
use chip_io_ovt_connects_horiz  gpio6_0_connects
timestamp 1706150479
transform -1 0 40840 0 -1 673770
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio6_0_pad
timestamp 1726580063
transform 0 -1 40000 1 0 645000
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio6_1_connects
timestamp 1706150479
transform -1 0 40840 0 -1 640770
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio6_1_pad
timestamp 1726580063
transform 0 -1 40000 1 0 612000
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio6_2_connects
timestamp 1706150479
transform -1 0 40840 0 -1 607770
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio6_2_pad
timestamp 1726580063
transform 0 -1 40000 1 0 579000
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio6_3_connects
timestamp 1706150479
transform -1 0 40840 0 -1 574770
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio6_3_pad
timestamp 1726580063
transform 0 -1 40000 1 0 546000
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio6_4_connects
timestamp 1706150479
transform -1 0 40840 0 -1 477170
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio6_4_pad
timestamp 1726580063
transform 0 -1 40000 1 0 448400
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio6_5_connects
timestamp 1706150479
transform -1 0 40840 0 -1 444170
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio6_5_pad
timestamp 1726580063
transform 0 -1 40000 1 0 415400
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio6_6_connects
timestamp 1706150479
transform -1 0 40840 0 -1 411170
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio6_6_pad
timestamp 1726580063
transform 0 -1 40000 1 0 382400
box -80 -147 28211 40151
use chip_io_ovt_connects_horiz  gpio6_7_connects
timestamp 1706150479
transform -1 0 40840 0 -1 378170
box 240 -2430 10095 28882
use sky130_fd_io__top_gpio_ovtv2  gpio6_7_pad
timestamp 1726580063
transform 0 -1 40000 1 0 349400
box -80 -147 28211 40151
use chip_io_gpio_connects_horiz  gpio7_0_connects
timestamp 1706150479
transform -1 0 40842 0 -1 282170
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio7_0_pad
timestamp 1726580063
transform 0 -1 39593 1 0 265400
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio7_1_connects
timestamp 1706150479
transform -1 0 40842 0 -1 261170
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio7_1_pad
timestamp 1726580063
transform 0 -1 39593 1 0 244400
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio7_2_connects
timestamp 1706150479
transform -1 0 40842 0 -1 240170
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio7_2_pad
timestamp 1726580063
transform 0 -1 39593 1 0 223400
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio7_3_connects
timestamp 1706150479
transform -1 0 40842 0 -1 219170
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio7_3_pad
timestamp 1726580063
transform 0 -1 39593 1 0 202400
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio7_4_connects
timestamp 1706150479
transform -1 0 40842 0 -1 155170
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio7_4_pad
timestamp 1726580063
transform 0 -1 39593 1 0 138400
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio7_5_connects
timestamp 1706150479
transform -1 0 40842 0 -1 134170
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio7_5_pad
timestamp 1726580063
transform 0 -1 39593 1 0 117400
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio7_6_connects
timestamp 1706150479
transform -1 0 40842 0 -1 113170
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio7_6_pad
timestamp 1726580063
transform 0 -1 39593 1 0 96400
box -143 -407 16134 39593
use chip_io_gpio_connects_horiz  gpio7_7_connects
timestamp 1706150479
transform -1 0 40842 0 -1 92170
box 0 -2430 10095 16814
use sky130_ef_io__gpiov2_pad  gpio7_7_pad
timestamp 1726580063
transform 0 -1 39593 1 0 75400
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio8_0_connects
timestamp 1726510233
transform 0 1 113343 -1 0 40910
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio8_0_pad
timestamp 1726580063
transform -1 0 130000 0 -1 39593
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio8_1_connects
timestamp 1726510233
transform 0 1 136343 -1 0 40910
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio8_1_pad
timestamp 1726580063
transform -1 0 153000 0 -1 39593
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio8_2_connects
timestamp 1726510233
transform 0 1 159343 -1 0 40910
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio8_2_pad
timestamp 1726580063
transform -1 0 176000 0 -1 39593
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio8_3_connects
timestamp 1726510233
transform 0 1 182343 -1 0 40910
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio8_3_pad
timestamp 1726580063
transform -1 0 199000 0 -1 39593
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio8_4_connects
timestamp 1726510233
transform 0 1 385343 -1 0 40910
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio8_4_pad
timestamp 1726580063
transform -1 0 402000 0 -1 39593
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio8_5_connects
timestamp 1726510233
transform 0 1 408343 -1 0 40910
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio8_5_pad
timestamp 1726580063
transform -1 0 425000 0 -1 39593
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio8_6_connects
timestamp 1726510233
transform 0 1 431343 -1 0 40910
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio8_6_pad
timestamp 1726580063
transform -1 0 448000 0 -1 39593
box -143 -407 16134 39593
use chip_io_gpio_connects_vert  gpio8_7_connects
timestamp 1726510233
transform 0 1 454343 -1 0 40910
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  gpio8_7_pad
timestamp 1726580063
transform -1 0 471000 0 -1 39593
box -143 -407 16134 39593
use muxsplit_connects  muxsplit_connects_ne
timestamp 1719074309
transform -1 0 677600 0 -1 996800
box 0 1305 300 7217
use muxsplit_connects  muxsplit_connects_nw
timestamp 1719074309
transform 1 0 40000 0 1 988000
box 0 1305 300 7217
use muxsplit_connects  muxsplit_connects_se
timestamp 1719074309
transform -1 0 677600 0 -1 49600
box 0 1305 300 7217
use muxsplit_connects  muxsplit_connects_sw
timestamp 1719074309
transform 1 0 40000 0 1 40800
box 0 1305 300 7217
use sky130_fd_io__top_amuxsplitv2  muxsplit_ne $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 0 1 677600 -1 0 996800
box 0 0 9600 40001
use sky130_fd_io__top_amuxsplitv2  muxsplit_nw
timestamp 1726580063
transform 0 -1 40000 1 0 988000
box 0 0 9600 40001
use sky130_fd_io__top_amuxsplitv2  muxsplit_se
timestamp 1726580063
transform 0 1 677600 -1 0 49600
box 0 0 9600 40001
use sky130_fd_io__top_amuxsplitv2  muxsplit_sw
timestamp 1726580063
transform 0 -1 40000 1 0 40800
box 0 0 9600 40001
use amuxbus_tap  n_amuxbus_tap
timestamp 1725852642
transform -1 0 369376 0 1 996600
box 0 0 1738 12222
use open_source  open_source_0
timestamp 1666123577
transform 1 0 675528 0 1 1013176
box 752 5164 29030 16242
use ovt_vinref_connects  ovt_vinref_connects_0
timestamp 1563079390
transform 1 0 0 0 1 0
box 39927 374670 677623 644952
use sky130_fd_io__top_pwrdetv2  pwrdet_s $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform -1 0 526180 0 -1 40000
box 282 0 10856 40000
use pwrdetv2_overlay  pwrdetv2_overlay_0
timestamp 1726600167
transform 1 0 8 0 1 2
box 518284 26330 524560 38196
use sky130_fd_io__top_xres4v2  resetb_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform -1 0 107000 0 -1 40000
box -103 0 15124 40000
use chip_io_gpio_connects_vert  select_connects
timestamp 1726510233
transform 0 1 68343 -1 0 40910
box 0 -2202 10158 16680
use sky130_ef_io__gpiov2_pad  select_pad
timestamp 1726580063
transform -1 0 85000 0 -1 39593
box -143 -407 16134 39593
use sky130_fd_io__top_sio_macro  sio_macro_pads $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform -1 0 670000 0 -1 50743
box 0 0 96000 50947
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform -1 0 676200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_1
timestamp 1726580063
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_2
timestamp 1726580063
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_3
timestamp 1726580063
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_4
timestamp 1726580063
transform 0 1 678007 -1 0 518200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_5
timestamp 1726580063
transform 1 0 676800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_6
timestamp 1726580063
transform 1 0 677000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_7
timestamp 1726580063
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_8
timestamp 1726580063
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  sky130_ef_io__com_bus_slice_1um_9
timestamp 1726580063
transform 0 -1 39593 1 0 520800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_1
timestamp 1726580063
transform -1 0 69000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_2
timestamp 1726580063
transform -1 0 92000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_3
timestamp 1726580063
transform -1 0 114000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_4
timestamp 1726580063
transform -1 0 137000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_5
timestamp 1726580063
transform -1 0 160000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_6
timestamp 1726580063
transform -1 0 183000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_7
timestamp 1726580063
transform -1 0 206000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_8
timestamp 1726580063
transform -1 0 228000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_9
timestamp 1726580063
transform -1 0 250000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_10
timestamp 1726580063
transform -1 0 272000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_11
timestamp 1726580063
transform -1 0 294000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_12
timestamp 1726580063
transform -1 0 316000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_13
timestamp 1726580063
transform -1 0 338000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_14
timestamp 1726580063
transform -1 0 360000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_15
timestamp 1726580063
transform -1 0 386000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_16
timestamp 1726580063
transform -1 0 409000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_17
timestamp 1726580063
transform -1 0 432000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_18
timestamp 1726580063
transform -1 0 455000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_19
timestamp 1726580063
transform -1 0 478000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_20
timestamp 1726580063
transform -1 0 500000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_21
timestamp 1726580063
transform -1 0 522000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_22
timestamp 1726580063
transform -1 0 548000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_23
timestamp 1726580063
transform -1 0 574000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_25
timestamp 1726580063
transform 0 1 678007 -1 0 74600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_26
timestamp 1726580063
transform 0 1 678007 -1 0 95600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_27
timestamp 1726580063
transform 0 1 678007 -1 0 116600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_28
timestamp 1726580063
transform 0 1 678007 -1 0 137600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_29
timestamp 1726580063
transform 0 1 678007 -1 0 158600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_30
timestamp 1726580063
transform 0 1 678007 -1 0 178600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_31
timestamp 1726580063
transform 0 1 678007 -1 0 198600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_32
timestamp 1726580063
transform 0 1 678007 -1 0 219600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_33
timestamp 1726580063
transform 0 1 678007 -1 0 240600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_34
timestamp 1726580063
transform 0 1 678007 -1 0 261600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_35
timestamp 1726580063
transform 0 1 678007 -1 0 282600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_36
timestamp 1726580063
transform 0 1 678007 -1 0 302600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_37
timestamp 1726580063
transform 0 1 678007 -1 0 322600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_38
timestamp 1726580063
transform 0 1 678007 -1 0 346600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_39
timestamp 1726580063
transform 0 1 678007 -1 0 379600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_40
timestamp 1726580063
transform 0 1 678007 -1 0 412600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_41
timestamp 1726580063
transform 0 1 678007 -1 0 445600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_42
timestamp 1726580063
transform 0 1 678007 -1 0 478600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_43
timestamp 1726580063
transform 0 1 678007 -1 0 498600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_44
timestamp 1726580063
transform 0 1 678007 -1 0 523200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_45
timestamp 1726580063
transform 0 1 678007 -1 0 543200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_46
timestamp 1726580063
transform 0 1 678007 -1 0 576200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_47
timestamp 1726580063
transform 0 1 678007 -1 0 609200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_48
timestamp 1726580063
transform 0 1 678007 -1 0 642200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_49
timestamp 1726580063
transform 0 1 678007 -1 0 675200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_50
timestamp 1726580063
transform 0 1 678007 -1 0 695200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_51
timestamp 1726580063
transform 0 1 678007 -1 0 715200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_52
timestamp 1726580063
transform 0 1 678007 -1 0 739200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_53
timestamp 1726580063
transform 0 1 678007 -1 0 759200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_54
timestamp 1726580063
transform 0 1 678007 -1 0 780200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_55
timestamp 1726580063
transform 0 1 678007 -1 0 801200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_56
timestamp 1726580063
transform 0 1 678007 -1 0 822200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_57
timestamp 1726580063
transform 0 1 678007 -1 0 843200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_58
timestamp 1726580063
transform 0 1 678007 -1 0 863200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_59
timestamp 1726580063
transform 0 1 678007 -1 0 884200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_60
timestamp 1726580063
transform 0 1 678007 -1 0 905200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_61
timestamp 1726580063
transform 0 1 678007 -1 0 926200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_62
timestamp 1726580063
transform 0 1 678007 -1 0 947200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_63
timestamp 1726580063
transform 0 1 678007 -1 0 967200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_64
timestamp 1726580063
transform 1 0 675800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_66
timestamp 1726580063
transform 0 -1 39593 1 0 74400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_67
timestamp 1726580063
transform 0 -1 39593 1 0 95400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_68
timestamp 1726580063
transform 0 -1 39593 1 0 116400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_69
timestamp 1726580063
transform 0 -1 39593 1 0 137400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_70
timestamp 1726580063
transform 0 -1 39593 1 0 158400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_71
timestamp 1726580063
transform 0 -1 39593 1 0 178400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_72
timestamp 1726580063
transform 0 -1 39593 1 0 181400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_73
timestamp 1726580063
transform 0 -1 39593 1 0 201400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_74
timestamp 1726580063
transform 0 -1 39593 1 0 222400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_75
timestamp 1726580063
transform 0 -1 39593 1 0 243400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_76
timestamp 1726580063
transform 0 -1 39593 1 0 264400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_77
timestamp 1726580063
transform 0 -1 39593 1 0 285400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_78
timestamp 1726580063
transform 0 -1 39593 1 0 305400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_79
timestamp 1726580063
transform 0 -1 39593 1 0 325400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_80
timestamp 1726580063
transform 0 -1 39593 1 0 328400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_81
timestamp 1726580063
transform 0 -1 39593 1 0 348400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_82
timestamp 1726580063
transform 0 -1 39593 1 0 381400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_83
timestamp 1726580063
transform 0 -1 39593 1 0 414400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_84
timestamp 1726580063
transform 0 -1 39593 1 0 447400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_85
timestamp 1726580063
transform 0 -1 39593 1 0 480400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_86
timestamp 1726580063
transform 0 -1 39593 1 0 500400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_87
timestamp 1726580063
transform 0 -1 39593 1 0 525000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_88
timestamp 1726580063
transform 0 -1 39593 1 0 545000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_89
timestamp 1726580063
transform 0 -1 39593 1 0 578000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_90
timestamp 1726580063
transform 0 -1 39593 1 0 611000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_91
timestamp 1726580063
transform 0 -1 39593 1 0 644000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_92
timestamp 1726580063
transform 0 -1 39593 1 0 677000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_93
timestamp 1726580063
transform 0 -1 39593 1 0 697000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_94
timestamp 1726580063
transform 0 -1 39593 1 0 717000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_95
timestamp 1726580063
transform 0 -1 39593 1 0 720000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_96
timestamp 1726580063
transform 0 -1 39593 1 0 740000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_97
timestamp 1726580063
transform 0 -1 39593 1 0 760000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_98
timestamp 1726580063
transform 0 -1 39593 1 0 781000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_99
timestamp 1726580063
transform 0 -1 39593 1 0 802000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_100
timestamp 1726580063
transform 0 -1 39593 1 0 823000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_101
timestamp 1726580063
transform 0 -1 39593 1 0 844000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_102
timestamp 1726580063
transform 0 -1 39593 1 0 864000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_103
timestamp 1726580063
transform 0 -1 39593 1 0 885000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_104
timestamp 1726580063
transform 0 -1 39593 1 0 906000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_105
timestamp 1726580063
transform 0 -1 39593 1 0 927000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_106
timestamp 1726580063
transform 0 -1 39593 1 0 948000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_107
timestamp 1726580063
transform 0 -1 39593 1 0 968000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  sky130_ef_io__com_bus_slice_5um_108
timestamp 1726580063
transform 0 -1 39593 1 0 971000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_1
timestamp 1726580063
transform -1 0 68000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_2
timestamp 1726580063
transform -1 0 91000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_3
timestamp 1726580063
transform -1 0 113000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_4
timestamp 1726580063
transform -1 0 136000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_5
timestamp 1726580063
transform -1 0 159000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_6
timestamp 1726580063
transform -1 0 182000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_7
timestamp 1726580063
transform -1 0 205000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_8
timestamp 1726580063
transform -1 0 227000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_9
timestamp 1726580063
transform -1 0 249000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_10
timestamp 1726580063
transform -1 0 271000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_11
timestamp 1726580063
transform -1 0 293000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_12
timestamp 1726580063
transform -1 0 315000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_13
timestamp 1726580063
transform -1 0 337000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_14
timestamp 1726580063
transform -1 0 359000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_15
timestamp 1726580063
transform -1 0 385000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_16
timestamp 1726580063
transform -1 0 408000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_17
timestamp 1726580063
transform -1 0 431000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_18
timestamp 1726580063
transform -1 0 454000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_19
timestamp 1726580063
transform -1 0 477000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_20
timestamp 1726580063
transform -1 0 499000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_21
timestamp 1726580063
transform -1 0 521000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_22
timestamp 1726580063
transform -1 0 547000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_23
timestamp 1726580063
transform -1 0 573000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_24
timestamp 1726580063
transform -1 0 676000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_25
timestamp 1726580063
transform 1 0 673800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_26
timestamp 1726580063
transform 0 -1 39593 1 0 179400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_27
timestamp 1726580063
transform 0 -1 39593 1 0 326400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_28
timestamp 1726580063
transform 0 -1 39593 1 0 718000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_10um  sky130_ef_io__com_bus_slice_10um_29
timestamp 1726580063
transform 0 -1 39593 1 0 969000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_1
timestamp 1726580063
transform -1 0 66000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_2
timestamp 1726580063
transform -1 0 89000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_3
timestamp 1726580063
transform -1 0 111000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_4
timestamp 1726580063
transform -1 0 134000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_5
timestamp 1726580063
transform -1 0 157000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_6
timestamp 1726580063
transform -1 0 180000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_7
timestamp 1726580063
transform -1 0 203000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_8
timestamp 1726580063
transform -1 0 225000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_9
timestamp 1726580063
transform -1 0 247000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_10
timestamp 1726580063
transform -1 0 269000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_11
timestamp 1726580063
transform -1 0 291000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_12
timestamp 1726580063
transform -1 0 313000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_13
timestamp 1726580063
transform -1 0 335000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_14
timestamp 1726580063
transform -1 0 357000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_15
timestamp 1726580063
transform -1 0 364000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_16
timestamp 1726580063
transform -1 0 383000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_17
timestamp 1726580063
transform -1 0 406000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_18
timestamp 1726580063
transform -1 0 429000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_19
timestamp 1726580063
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_20
timestamp 1726580063
transform -1 0 475000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_21
timestamp 1726580063
transform -1 0 497000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_22
timestamp 1726580063
transform -1 0 519000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_23
timestamp 1726580063
transform -1 0 526000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_24
timestamp 1726580063
transform -1 0 545000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_25
timestamp 1726580063
transform -1 0 571000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_26
timestamp 1726580063
transform -1 0 674000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_27
timestamp 1726580063
transform 0 1 678007 -1 0 53600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_28
timestamp 1726580063
transform 0 1 678007 -1 0 73600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_29
timestamp 1726580063
transform 0 1 678007 -1 0 94600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_30
timestamp 1726580063
transform 0 1 678007 -1 0 115600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_31
timestamp 1726580063
transform 0 1 678007 -1 0 136600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_32
timestamp 1726580063
transform 0 1 678007 -1 0 157600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_33
timestamp 1726580063
transform 0 1 678007 -1 0 177600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_34
timestamp 1726580063
transform 0 1 678007 -1 0 197600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_35
timestamp 1726580063
transform 0 1 678007 -1 0 218600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_36
timestamp 1726580063
transform 0 1 678007 -1 0 239600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_37
timestamp 1726580063
transform 0 1 678007 -1 0 260600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_38
timestamp 1726580063
transform 0 1 678007 -1 0 281600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_39
timestamp 1726580063
transform 0 1 678007 -1 0 301600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_40
timestamp 1726580063
transform 0 1 678007 -1 0 321600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_41
timestamp 1726580063
transform 0 1 678007 -1 0 326600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_42
timestamp 1726580063
transform 0 1 678007 -1 0 345600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_43
timestamp 1726580063
transform 0 1 678007 -1 0 378600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_44
timestamp 1726580063
transform 0 1 678007 -1 0 411600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_45
timestamp 1726580063
transform 0 1 678007 -1 0 444600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_46
timestamp 1726580063
transform 0 1 678007 -1 0 477600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_47
timestamp 1726580063
transform 0 1 678007 -1 0 497600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_48
timestamp 1726580063
transform 0 1 678007 -1 0 522200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_49
timestamp 1726580063
transform 0 1 678007 -1 0 542200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_50
timestamp 1726580063
transform 0 1 678007 -1 0 575200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_51
timestamp 1726580063
transform 0 1 678007 -1 0 608200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_52
timestamp 1726580063
transform 0 1 678007 -1 0 641200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_53
timestamp 1726580063
transform 0 1 678007 -1 0 674200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_54
timestamp 1726580063
transform 0 1 678007 -1 0 694200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_55
timestamp 1726580063
transform 0 1 678007 -1 0 714200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_56
timestamp 1726580063
transform 0 1 678007 -1 0 719200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_57
timestamp 1726580063
transform 0 1 678007 -1 0 738200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_58
timestamp 1726580063
transform 0 1 678007 -1 0 758200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_59
timestamp 1726580063
transform 0 1 678007 -1 0 779200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_60
timestamp 1726580063
transform 0 1 678007 -1 0 800200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_61
timestamp 1726580063
transform 0 1 678007 -1 0 821200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_62
timestamp 1726580063
transform 0 1 678007 -1 0 842200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_63
timestamp 1726580063
transform 0 1 678007 -1 0 862200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_64
timestamp 1726580063
transform 0 1 678007 -1 0 883200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_65
timestamp 1726580063
transform 0 1 678007 -1 0 904200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_66
timestamp 1726580063
transform 0 1 678007 -1 0 925200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_67
timestamp 1726580063
transform 0 1 678007 -1 0 946200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_68
timestamp 1726580063
transform 0 1 678007 -1 0 966200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_69
timestamp 1726580063
transform 0 1 678007 -1 0 971200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_70
timestamp 1726580063
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_71
timestamp 1726580063
transform 1 0 59800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_72
timestamp 1726580063
transform 1 0 63800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_73
timestamp 1726580063
transform 1 0 83800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_74
timestamp 1726580063
transform 1 0 87800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_75
timestamp 1726580063
transform 1 0 107800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_76
timestamp 1726580063
transform 1 0 111800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_77
timestamp 1726580063
transform 1 0 131800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_78
timestamp 1726580063
transform 1 0 135800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_79
timestamp 1726580063
transform 1 0 155800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_80
timestamp 1726580063
transform 1 0 159800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_81
timestamp 1726580063
transform 1 0 178800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_82
timestamp 1726580063
transform 1 0 182800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_83
timestamp 1726580063
transform 1 0 201800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_84
timestamp 1726580063
transform 1 0 205800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_85
timestamp 1726580063
transform 1 0 225800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_86
timestamp 1726580063
transform 1 0 229800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_87
timestamp 1726580063
transform 1 0 249800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_88
timestamp 1726580063
transform 1 0 253800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_89
timestamp 1726580063
transform 1 0 273800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_90
timestamp 1726580063
transform 1 0 277800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_91
timestamp 1726580063
transform 1 0 297800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_92
timestamp 1726580063
transform 1 0 301800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_93
timestamp 1726580063
transform 1 0 320800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_94
timestamp 1726580063
transform 1 0 324800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_95
timestamp 1726580063
transform 1 0 343800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_96
timestamp 1726580063
transform 1 0 347800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_97
timestamp 1726580063
transform 1 0 366800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_98
timestamp 1726580063
transform 1 0 370800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_99
timestamp 1726580063
transform 1 0 389800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_100
timestamp 1726580063
transform 1 0 393800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_101
timestamp 1726580063
transform 1 0 412800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_102
timestamp 1726580063
transform 1 0 416800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_103
timestamp 1726580063
transform 1 0 436800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_104
timestamp 1726580063
transform 1 0 440800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_105
timestamp 1726580063
transform 1 0 460800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_106
timestamp 1726580063
transform 1 0 464800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_107
timestamp 1726580063
transform 1 0 484800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_108
timestamp 1726580063
transform 1 0 488800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_109
timestamp 1726580063
transform 1 0 508800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_110
timestamp 1726580063
transform 1 0 512800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_111
timestamp 1726580063
transform 1 0 531800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_112
timestamp 1726580063
transform 1 0 535800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_113
timestamp 1726580063
transform 1 0 554800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_114
timestamp 1726580063
transform 1 0 558800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_115
timestamp 1726580063
transform 1 0 578800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_116
timestamp 1726580063
transform 1 0 582800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_117
timestamp 1726580063
transform 1 0 602800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_118
timestamp 1726580063
transform 1 0 606800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_119
timestamp 1726580063
transform 1 0 626800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_120
timestamp 1726580063
transform 1 0 630800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_121
timestamp 1726580063
transform 1 0 650800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_122
timestamp 1726580063
transform 1 0 654800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_123
timestamp 1726580063
transform 0 -1 39593 1 0 50400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_124
timestamp 1726580063
transform 0 -1 39593 1 0 70400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_125
timestamp 1726580063
transform 0 -1 39593 1 0 91400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_126
timestamp 1726580063
transform 0 -1 39593 1 0 112400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_127
timestamp 1726580063
transform 0 -1 39593 1 0 133400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_128
timestamp 1726580063
transform 0 -1 39593 1 0 154400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_129
timestamp 1726580063
transform 0 -1 39593 1 0 174400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_130
timestamp 1726580063
transform 0 -1 39593 1 0 197400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_131
timestamp 1726580063
transform 0 -1 39593 1 0 218400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_132
timestamp 1726580063
transform 0 -1 39593 1 0 239400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_133
timestamp 1726580063
transform 0 -1 39593 1 0 260400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_134
timestamp 1726580063
transform 0 -1 39593 1 0 281400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_135
timestamp 1726580063
transform 0 -1 39593 1 0 301400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_136
timestamp 1726580063
transform 0 -1 39593 1 0 321400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_137
timestamp 1726580063
transform 0 -1 39593 1 0 344400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_138
timestamp 1726580063
transform 0 -1 39593 1 0 377400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_139
timestamp 1726580063
transform 0 -1 39593 1 0 410400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_140
timestamp 1726580063
transform 0 -1 39593 1 0 443400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_141
timestamp 1726580063
transform 0 -1 39593 1 0 476400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_142
timestamp 1726580063
transform 0 -1 39593 1 0 496400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_143
timestamp 1726580063
transform 0 -1 39593 1 0 521000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_144
timestamp 1726580063
transform 0 -1 39593 1 0 541000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_145
timestamp 1726580063
transform 0 -1 39593 1 0 574000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_146
timestamp 1726580063
transform 0 -1 39593 1 0 607000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_147
timestamp 1726580063
transform 0 -1 39593 1 0 640000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_148
timestamp 1726580063
transform 0 -1 39593 1 0 673000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_149
timestamp 1726580063
transform 0 -1 39593 1 0 693000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_150
timestamp 1726580063
transform 0 -1 39593 1 0 713000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_151
timestamp 1726580063
transform 0 -1 39593 1 0 736000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_152
timestamp 1726580063
transform 0 -1 39593 1 0 756000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_153
timestamp 1726580063
transform 0 -1 39593 1 0 777000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_154
timestamp 1726580063
transform 0 -1 39593 1 0 798000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_155
timestamp 1726580063
transform 0 -1 39593 1 0 819000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_156
timestamp 1726580063
transform 0 -1 39593 1 0 840000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_157
timestamp 1726580063
transform 0 -1 39593 1 0 860000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_158
timestamp 1726580063
transform 0 -1 39593 1 0 881000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_159
timestamp 1726580063
transform 0 -1 39593 1 0 902000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_160
timestamp 1726580063
transform 0 -1 39593 1 0 923000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_161
timestamp 1726580063
transform 0 -1 39593 1 0 944000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  sky130_ef_io__com_bus_slice_20um_162
timestamp 1726580063
transform 0 -1 39593 1 0 964000
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform -1 0 552000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  sky130_ef_io__disconnect_vdda_slice_5um_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 0 1 678007 -1 0 987200
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  sky130_ef_io__disconnect_vdda_slice_5um_1
timestamp 1726580063
transform 0 -1 39593 1 0 987000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  sky130_ef_io__disconnect_vdda_slice_5um_2
timestamp 1726580063
transform 0 -1 39593 1 0 54400
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  sky130_ef_io__disconnect_vdda_slice_5um_3
timestamp 1726580063
transform 0 1 678007 -1 0 54600
box 0 0 1000 39593
use user_id_textblock  user_id_textblock_0
timestamp 1608324878
transform 1 0 12306 0 1 9642
box -656 1508 33720 10344
use sky130_fd_io__top_vrefcapv2  vcap_e $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 0 1 677600 -1 0 518056
box 0 0 3456 40000
use sky130_fd_io__top_vrefcapv2  vcap_w
timestamp 1726580063
transform 0 -1 40000 1 0 517400
box 0 0 3456 40000
use sky130_ef_io__vccd_lvc_clamped_pad  vccd0_0_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform -1 0 62000 0 -1 39593
box 0 -2107 17239 39593
use sky130_ef_io__vccd_lvc_clamped_pad  vccd0_1_pad
timestamp 1726580063
transform -1 0 379000 0 -1 39593
box 0 -2107 17239 39593
use sky130_ef_io__vccd_lvc_clamped3_pad  vccd1_0_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 0 1 678007 -1 0 493600
box 0 -2177 17187 39593
use sky130_ef_io__vccd_lvc_clamped3_pad  vccd1_1_pad
timestamp 1726580063
transform 0 1 678007 -1 0 962200
box 0 -2177 17187 39593
use sky130_ef_io__vccd_lvc_clamped3_pad  vccd1_2_pad
timestamp 1726580063
transform 1 0 516800 0 1 998007
box 0 -2177 17187 39593
use sky130_ef_io__vccd_lvc_clamped3_pad  vccd2_0_pad
timestamp 1726580063
transform 1 0 44800 0 1 998007
box 0 -2177 17187 39593
use sky130_ef_io__vccd_lvc_clamped3_pad  vccd2_1_pad
timestamp 1726580063
transform 0 -1 39593 1 0 741000
box 0 -2177 17187 39593
use sky130_ef_io__vccd_lvc_clamped3_pad  vccd2_2_pad
timestamp 1726580063
transform 0 -1 39593 1 0 159400
box 0 -2177 17187 39593
use sky130_ef_io__vdda_hvc_clamped_pad  vdda0_0_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 1 0 374800 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  vdda1_0_pad
timestamp 1726580063
transform 0 1 678007 -1 0 317600
box 0 -407 15000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  vdda1_1_pad
timestamp 1726580063
transform 0 1 678007 -1 0 710200
box 0 -407 15000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  vdda2_0_pad
timestamp 1726580063
transform 0 -1 39593 1 0 698000
box 0 -407 15000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  vdda2_1_pad
timestamp 1726580063
transform 0 -1 39593 1 0 306400
box 0 -407 15000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  vdda3_0_pad
timestamp 1726580063
transform -1 0 541000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  vddio_0_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 0 1 678007 -1 0 69600
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  vddio_1_pad
timestamp 1726580063
transform 0 1 678007 -1 0 297600
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  vddio_2_pad
timestamp 1726580063
transform 0 1 678007 -1 0 690200
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  vddio_3_pad
timestamp 1726580063
transform 0 1 678007 -1 0 986200
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  vddio_4_pad
timestamp 1726580063
transform 1 0 397800 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  vddio_5_pad
timestamp 1726580063
transform 0 -1 39593 1 0 972000
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  vddio_6_pad
timestamp 1726580063
transform 0 -1 39593 1 0 678000
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  vddio_7_pad
timestamp 1726580063
transform 0 -1 39593 1 0 286400
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  vddio_8_pad
timestamp 1726580063
transform 0 -1 39593 1 0 55400
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  vddio_9_pad
timestamp 1726580063
transform -1 0 353000 0 -1 39593
box 0 -407 15000 39593
use vref_connects  vref_connects_e
timestamp 1726510490
transform -1 0 677600 0 -1 514600
box 0 972 300 13139
use vref_connects  vref_connects_w
timestamp 1726510490
transform 1 0 40000 0 1 501400
box 0 972 300 13139
use sky130_fd_io__top_gpiovrefv2  vref_e $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 0 1 677600 -1 0 514600
box 0 0 16000 40000
use sky130_fd_io__top_gpiovrefv2  vref_w
timestamp 1726580063
transform 0 -1 40000 1 0 501400
box 0 0 16000 40000
use sky130_ef_io__vssa_hvc_clamped_pad  vssa0_0_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 1 0 305800 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  vssa1_0_pad
timestamp 1726580063
transform 0 1 678007 -1 0 341600
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  vssa1_1_pad
timestamp 1726580063
transform 0 1 678007 -1 0 734200
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  vssa2_0_pad
timestamp 1726580063
transform 0 -1 39593 1 0 721000
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  vssa2_1_pad
timestamp 1726580063
transform 0 -1 39593 1 0 329400
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  vssa3_0_pad
timestamp 1726580063
transform -1 0 515000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped_pad  vssd0_0_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform -1 0 243000 0 -1 39593
box 0 -2107 17239 39593
use sky130_ef_io__vssd_lvc_clamped_pad  vssd0_1_pad
timestamp 1726580063
transform -1 0 567000 0 -1 39593
box 0 -2107 17239 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  vssd1_0_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 0 1 678007 -1 0 173600
box 0 -2177 17187 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  vssd1_1_pad
timestamp 1726580063
transform 0 1 678007 -1 0 754200
box 0 -2177 17187 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  vssd1_2_pad
timestamp 1726580063
transform 1 0 658800 0 1 998007
box 0 -2177 17187 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  vssd2_0_pad
timestamp 1726580063
transform 1 0 186800 0 1 998007
box 0 -2177 17187 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  vssd2_1_pad
timestamp 1726580063
transform 0 -1 39593 1 0 949000
box 0 -2177 17187 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  vssd2_2_pad
timestamp 1726580063
transform 0 -1 39593 1 0 481400
box 0 -2177 17187 39593
use sky130_ef_io__vssio_hvc_clamped_pad  vssio_0_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1726580063
transform 0 1 678007 -1 0 193600
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  vssio_1_pad
timestamp 1726580063
transform 0 1 678007 -1 0 538200
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  vssio_2_pad
timestamp 1726580063
transform 0 1 678007 -1 0 858200
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  vssio_3_pad
timestamp 1726580063
transform 1 0 539800 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  vssio_4_pad
timestamp 1726580063
transform 1 0 163800 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  vssio_5_pad
timestamp 1726580063
transform 0 -1 39593 1 0 845000
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  vssio_6_pad
timestamp 1726580063
transform 0 -1 39593 1 0 526000
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  vssio_7_pad
timestamp 1726580063
transform 0 -1 39593 1 0 182400
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  vssio_8_pad
timestamp 1726580063
transform -1 0 221000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  vssio_9_pad
timestamp 1726580063
transform -1 0 493000 0 -1 39593
box 0 -407 15000 39593
use sky130_fd_io__top_analog_pad  xi0_pad
timestamp 1726580063
transform -1 0 265000 0 -1 39600
box -80 0 15080 39600
use sky130_fd_io__top_analog_pad  xi1_pad
timestamp 1726580063
transform -1 0 309000 0 -1 39600
box -80 0 15080 39600
use sky130_fd_io__top_analog_pad  xo0_pad
timestamp 1726580063
transform -1 0 287000 0 -1 39600
box -80 0 15080 39600
use sky130_fd_io__top_analog_pad  xo1_pad
timestamp 1726580063
transform -1 0 331000 0 -1 39600
box -80 0 15080 39600
<< labels >>
flabel metal5 s 50500 8920 58500 16920 0 FreeSans 24000 0 0 0 vccd0_0
port 1 nsew power bidirectional
flabel metal5 s 72500 8843 80500 16843 0 FreeSans 24000 0 0 0 select
port 2 nsew signal bidirectional
flabel metal5 s 95500 8920 103500 16920 0 FreeSans 24000 0 0 0 resetb
port 3 nsew signal input
flabel metal5 s 117500 8843 125500 16843 0 FreeSans 24000 0 0 0 gpio8_0
port 4 nsew signal bidirectional
flabel metal5 s 140500 8843 148500 16843 0 FreeSans 24000 0 0 0 gpio8_1
port 5 nsew signal bidirectional
flabel metal5 s 163500 8843 171500 16843 0 FreeSans 24000 0 0 0 gpio8_2
port 6 nsew signal bidirectional
flabel metal5 s 186500 8843 194500 16843 0 FreeSans 24000 0 0 0 gpio8_3
port 7 nsew signal bidirectional
flabel metal5 s 209500 8920 217500 16920 0 FreeSans 24000 0 0 0 vssio_8
port 8 nsew ground bidirectional
flabel metal5 s 231500 8920 239500 16920 0 FreeSans 24000 0 0 0 vssd0_0
port 9 nsew ground bidirectional
flabel metal5 s 253500 8920 261500 16920 0 FreeSans 24000 0 0 0 xi0
port 10 nsew signal bidirectional
flabel metal5 s 275500 8920 283500 16920 0 FreeSans 24000 0 0 0 xo0
port 11 nsew signal bidirectional
flabel metal5 s 297500 8920 305500 16920 0 FreeSans 24000 0 0 0 xi1
port 12 nsew signal bidirectional
flabel metal5 s 319500 8920 327500 16920 0 FreeSans 24000 0 0 0 xo1
port 13 nsew signal bidirectional
flabel metal5 s 341500 8920 349500 16920 0 FreeSans 24000 0 0 0 vddio_9
port 14 nsew power bidirectional
flabel metal5 s 367500 8920 375500 16920 0 FreeSans 24000 0 0 0 vccd0_1
port 15 nsew power bidirectional
flabel metal5 s 389500 8843 397500 16843 0 FreeSans 24000 0 0 0 gpio8_4
port 16 nsew signal bidirectional
flabel metal5 s 412500 8843 420500 16843 0 FreeSans 24000 0 0 0 gpio8_5
port 17 nsew signal bidirectional
flabel metal5 s 435500 8843 443500 16843 0 FreeSans 24000 0 0 0 gpio8_6
port 18 nsew signal bidirectional
flabel metal5 s 458500 8843 466500 16843 0 FreeSans 24000 0 0 0 gpio8_7
port 19 nsew signal bidirectional
flabel metal5 s 481500 8920 489500 16920 0 FreeSans 24000 0 0 0 vssio_9
port 20 nsew ground bidirectional
flabel metal5 s 503500 8920 511500 16920 0 FreeSans 24000 0 0 0 vssa3_0
port 21 nsew ground bidirectional
flabel metal5 s 529500 8920 537500 16920 0 FreeSans 24000 0 0 0 vdda3_0
port 22 nsew power bidirectional
flabel metal5 s 555500 8920 563500 16920 0 FreeSans 24000 0 0 0 vssd0_1
port 23 nsew ground bidirectional
flabel metal5 s 615697 14068 623697 22068 0 FreeSans 24000 0 0 0 sio0
port 24 nsew signal bidirectional
flabel metal5 s 638302 14068 646302 22068 0 FreeSans 24000 0 0 0 sio1
port 25 nsew signal bidirectional
flabel metal5 s 700680 58100 708680 66100 0 FreeSans 24000 0 0 0 vddio_0
port 26 nsew power bidirectional
flabel metal5 s 700757 78100 708757 86100 0 FreeSans 24000 0 0 0 gpio0_0
port 27 nsew signal bidirectional
flabel metal5 s 700757 99100 708757 107100 0 FreeSans 24000 0 0 0 gpio0_1
port 28 nsew signal bidirectional
flabel metal5 s 700757 120100 708757 128100 0 FreeSans 24000 0 0 0 gpio0_2
port 29 nsew signal bidirectional
flabel metal5 s 700757 141100 708757 149100 0 FreeSans 24000 0 0 0 gpio0_3
port 30 nsew signal bidirectional
flabel metal5 s 700680 162100 708680 170100 0 FreeSans 24000 0 0 0 vssd1_0
port 31 nsew ground bidirectional
flabel metal5 s 700680 182100 708680 190100 0 FreeSans 24000 0 0 0 vssio_0
port 32 nsew ground bidirectional
flabel metal5 s 700757 202100 708757 210100 0 FreeSans 24000 0 0 0 gpio0_4
port 33 nsew signal bidirectional
flabel metal5 s 700757 223100 708757 231100 0 FreeSans 24000 0 0 0 gpio0_5
port 34 nsew signal bidirectional
flabel metal5 s 700757 244100 708757 252100 0 FreeSans 24000 0 0 0 gpio0_6
port 35 nsew signal bidirectional
flabel metal5 s 700757 265100 708757 273100 0 FreeSans 24000 0 0 0 gpio0_7
port 36 nsew signal bidirectional
flabel metal5 s 700680 286100 708680 294100 0 FreeSans 24000 0 0 0 vddio_1
port 37 nsew power bidirectional
flabel metal5 s 700680 306100 708680 314100 0 FreeSans 24000 0 0 0 vdda1_0
port 38 nsew power bidirectional
flabel metal5 s 700680 330100 708680 338100 0 FreeSans 24000 0 0 0 vssa1_0
port 39 nsew ground bidirectional
flabel metal5 s 701096 359734 709096 367734 0 FreeSans 24000 0 0 0 gpio1_0
port 40 nsew signal bidirectional
flabel metal5 s 701096 392734 709096 400734 0 FreeSans 24000 0 0 0 gpio1_1
port 41 nsew signal bidirectional
flabel metal5 s 701096 425734 709096 433734 0 FreeSans 24000 0 0 0 gpio1_2
port 42 nsew signal bidirectional
flabel metal5 s 701096 458734 709096 466734 0 FreeSans 24000 0 0 0 gpio1_3
port 43 nsew signal bidirectional
flabel metal5 s 700680 482100 708680 490100 0 FreeSans 24000 0 0 0 vccd1_0
port 44 nsew power bidirectional
flabel metal5 s 700680 526700 708680 534700 0 FreeSans 24000 0 0 0 vssio_1
port 45 nsew ground bidirectional
flabel metal5 s 701096 556334 709096 564334 0 FreeSans 24000 0 0 0 gpio1_4
port 46 nsew signal bidirectional
flabel metal5 s 701096 589334 709096 597334 0 FreeSans 24000 0 0 0 gpio1_5
port 47 nsew signal bidirectional
flabel metal5 s 701096 622334 709096 630334 0 FreeSans 24000 0 0 0 gpio1_6
port 48 nsew signal bidirectional
flabel metal5 s 701096 655334 709096 663334 0 FreeSans 24000 0 0 0 gpio1_7
port 49 nsew signal bidirectional
flabel metal5 s 700680 678700 708680 686700 0 FreeSans 24000 0 0 0 vddio_2
port 50 nsew power bidirectional
flabel metal5 s 700680 698700 708680 706700 0 FreeSans 24000 0 0 0 vdda1_1
port 51 nsew power bidirectional
flabel metal5 s 700680 722700 708680 730700 0 FreeSans 24000 0 0 0 vssa1_1
port 52 nsew ground bidirectional
flabel metal5 s 700680 742700 708680 750700 0 FreeSans 24000 0 0 0 vssd1_1
port 53 nsew ground bidirectional
flabel metal5 s 700757 762700 708757 770700 0 FreeSans 24000 0 0 0 gpio2_0
port 54 nsew signal bidirectional
flabel metal5 s 700757 783700 708757 791700 0 FreeSans 24000 0 0 0 gpio2_1
port 55 nsew signal bidirectional
flabel metal5 s 700757 804700 708757 812700 0 FreeSans 24000 0 0 0 gpio2_2
port 56 nsew signal bidirectional
flabel metal5 s 700757 825700 708757 833700 0 FreeSans 24000 0 0 0 gpio2_3
port 57 nsew signal bidirectional
flabel metal5 s 700680 846700 708680 854700 0 FreeSans 24000 0 0 0 vssio_2
port 58 nsew ground bidirectional
flabel metal5 s 700757 866700 708757 874700 0 FreeSans 24000 0 0 0 gpio2_4
port 59 nsew signal bidirectional
flabel metal5 s 700757 887700 708757 895700 0 FreeSans 24000 0 0 0 gpio2_5
port 60 nsew signal bidirectional
flabel metal5 s 700757 908700 708757 916700 0 FreeSans 24000 0 0 0 gpio2_6
port 61 nsew signal bidirectional
flabel metal5 s 700757 929700 708757 937700 0 FreeSans 24000 0 0 0 gpio2_7
port 62 nsew signal bidirectional
flabel metal5 s 700680 950700 708680 958700 0 FreeSans 24000 0 0 0 vccd1_1
port 63 nsew power bidirectional
flabel metal5 s 700680 974700 708680 982700 0 FreeSans 24000 0 0 0 vddio_3
port 64 nsew power bidirectional
flabel metal5 s 48300 1020680 56300 1028680 0 FreeSans 24000 0 0 0 vccd2_0
port 65 nsew power bidirectional
flabel metal5 s 72300 1020757 80300 1028757 0 FreeSans 24000 0 0 0 gpio4_7
port 66 nsew signal bidirectional
flabel metal5 s 96300 1020757 104300 1028757 0 FreeSans 24000 0 0 0 gpio4_6
port 67 nsew signal bidirectional
flabel metal5 s 120300 1020757 128300 1028757 0 FreeSans 24000 0 0 0 gpio4_5
port 68 nsew signal bidirectional
flabel metal5 s 144300 1020757 152300 1028757 0 FreeSans 24000 0 0 0 gpio4_4
port 69 nsew signal bidirectional
flabel metal5 s 167300 1020680 175300 1028680 0 FreeSans 24000 0 0 0 vssio_4
port 70 nsew ground bidirectional
flabel metal5 s 190300 1020680 198300 1028680 0 FreeSans 24000 0 0 0 vssd2_0
port 71 nsew ground bidirectional
flabel metal5 s 214300 1020757 222300 1028757 0 FreeSans 24000 0 0 0 gpio4_3
port 72 nsew signal bidirectional
flabel metal5 s 238300 1020757 246300 1028757 0 FreeSans 24000 0 0 0 gpio4_2
port 73 nsew signal bidirectional
flabel metal5 s 262300 1020757 270300 1028757 0 FreeSans 24000 0 0 0 gpio4_1
port 74 nsew signal bidirectional
flabel metal5 s 286300 1020757 294300 1028757 0 FreeSans 24000 0 0 0 gpio4_0
port 75 nsew signal bidirectional
flabel metal5 s 309300 1020680 317300 1028680 0 FreeSans 24000 0 0 0 vssa0_0
port 76 nsew ground bidirectional
flabel metal5 s 332300 1020680 340300 1028680 0 FreeSans 24000 0 0 0 analog_1
port 77 nsew signal bidirectional
flabel metal5 s 355300 1020680 363300 1028680 0 FreeSans 24000 0 0 0 analog_0
port 78 nsew signal bidirectional
flabel metal5 s 378300 1020680 386300 1028680 0 FreeSans 24000 0 0 0 vdda0_0
port 79 nsew power bidirectional
flabel metal5 s 401300 1020680 409300 1028680 0 FreeSans 24000 0 0 0 vddio_4
port 80 nsew power bidirectional
flabel metal5 s 425300 1020757 433300 1028757 0 FreeSans 24000 0 0 0 gpio3_7
port 81 nsew signal bidirectional
flabel metal5 s 449300 1020757 457300 1028757 0 FreeSans 24000 0 0 0 gpio3_6
port 82 nsew signal bidirectional
flabel metal5 s 473300 1020757 481300 1028757 0 FreeSans 24000 0 0 0 gpio3_5
port 83 nsew signal bidirectional
flabel metal5 s 497300 1020757 505300 1028757 0 FreeSans 24000 0 0 0 gpio3_4
port 84 nsew signal bidirectional
flabel metal5 s 520300 1020680 528300 1028680 0 FreeSans 24000 0 0 0 vccd1_2
port 85 nsew power bidirectional
flabel metal5 s 543300 1020680 551300 1028680 0 FreeSans 24000 0 0 0 vssio_3
port 86 nsew ground bidirectional
flabel metal5 s 567300 1020757 575300 1028757 0 FreeSans 24000 0 0 0 gpio3_3
port 87 nsew signal bidirectional
flabel metal5 s 591300 1020757 599300 1028757 0 FreeSans 24000 0 0 0 gpio3_2
port 88 nsew signal bidirectional
flabel metal5 s 615300 1020757 623300 1028757 0 FreeSans 24000 0 0 0 gpio3_1
port 89 nsew signal bidirectional
flabel metal5 s 639300 1020757 647300 1028757 0 FreeSans 24000 0 0 0 gpio3_0
port 90 nsew signal bidirectional
flabel metal5 s 662300 1020680 670300 1028680 0 FreeSans 24000 0 0 0 vssd1_2
port 91 nsew ground bidirectional
flabel metal5 s 8920 58900 16920 66900 0 FreeSans 24000 0 0 0 vddio_8
port 92 nsew power bidirectional
flabel metal5 s 8843 79900 16843 87900 0 FreeSans 24000 0 0 0 gpio7_7
port 93 nsew signal bidirectional
flabel metal5 s 8843 100900 16843 108900 0 FreeSans 24000 0 0 0 gpio7_6
port 94 nsew signal bidirectional
flabel metal5 s 8843 121900 16843 129900 0 FreeSans 24000 0 0 0 gpio7_5
port 95 nsew signal bidirectional
flabel metal5 s 8843 142900 16843 150900 0 FreeSans 24000 0 0 0 gpio7_4
port 96 nsew signal bidirectional
flabel metal5 s 8920 162900 16920 170900 0 FreeSans 24000 0 0 0 vccd2_2
port 97 nsew power bidirectional
flabel metal5 s 8920 185900 16920 193900 0 FreeSans 24000 0 0 0 vssio_7
port 98 nsew ground bidirectional
flabel metal5 s 8843 206900 16843 214900 0 FreeSans 24000 0 0 0 gpio7_3
port 99 nsew signal bidirectional
flabel metal5 s 8843 227900 16843 235900 0 FreeSans 24000 0 0 0 gpio7_2
port 100 nsew signal bidirectional
flabel metal5 s 8843 248900 16843 256900 0 FreeSans 24000 0 0 0 gpio7_1
port 101 nsew signal bidirectional
flabel metal5 s 8843 269900 16843 277900 0 FreeSans 24000 0 0 0 gpio7_0
port 102 nsew signal bidirectional
flabel metal5 s 8920 289900 16920 297900 0 FreeSans 24000 0 0 0 vddio_7
port 103 nsew power bidirectional
flabel metal5 s 8920 309900 16920 317900 0 FreeSans 24000 0 0 0 vdda2_1
port 104 nsew power bidirectional
flabel metal5 s 8920 332900 16920 340900 0 FreeSans 24000 0 0 0 vssa2_1
port 105 nsew ground bidirectional
flabel metal5 s 8504 356266 16504 364266 0 FreeSans 24000 0 0 0 gpio6_7
port 106 nsew signal bidirectional
flabel metal5 s 8504 389266 16504 397266 0 FreeSans 24000 0 0 0 gpio6_6
port 107 nsew signal bidirectional
flabel metal5 s 8504 422266 16504 430266 0 FreeSans 24000 0 0 0 gpio6_5
port 108 nsew signal bidirectional
flabel metal5 s 8504 455266 16504 463266 0 FreeSans 24000 0 0 0 gpio6_4
port 109 nsew signal bidirectional
flabel metal5 s 8920 484900 16920 492900 0 FreeSans 24000 0 0 0 vssd2_2
port 110 nsew ground bidirectional
flabel metal5 s 8920 529500 16920 537500 0 FreeSans 24000 0 0 0 vssio_6
port 111 nsew ground bidirectional
flabel metal5 s 8504 552866 16504 560866 0 FreeSans 24000 0 0 0 gpio6_3
port 112 nsew signal bidirectional
flabel metal5 s 8504 585866 16504 593866 0 FreeSans 24000 0 0 0 gpio6_2
port 113 nsew signal bidirectional
flabel metal5 s 8504 618866 16504 626866 0 FreeSans 24000 0 0 0 gpio6_1
port 114 nsew signal bidirectional
flabel metal5 s 8504 651866 16504 659866 0 FreeSans 24000 0 0 0 gpio6_0
port 115 nsew signal bidirectional
flabel metal5 s 8920 681500 16920 689500 0 FreeSans 24000 0 0 0 vddio_6
port 116 nsew power bidirectional
flabel metal5 s 8920 701500 16920 709500 0 FreeSans 24000 0 0 0 vdda2_0
port 117 nsew power bidirectional
flabel metal5 s 8920 724500 16920 732500 0 FreeSans 24000 0 0 0 vssa2_0
port 118 nsew ground bidirectional
flabel metal5 s 8920 744500 16920 752500 0 FreeSans 24000 0 0 0 vccd2_1
port 119 nsew power bidirectional
flabel metal5 s 8843 765500 16843 773500 0 FreeSans 24000 0 0 0 gpio5_7
port 120 nsew signal bidirectional
flabel metal5 s 8843 786500 16843 794500 0 FreeSans 24000 0 0 0 gpio5_6
port 121 nsew signal bidirectional
flabel metal5 s 8843 807500 16843 815500 0 FreeSans 24000 0 0 0 gpio5_5
port 122 nsew signal bidirectional
flabel metal5 s 8843 828500 16843 836500 0 FreeSans 24000 0 0 0 gpio5_4
port 123 nsew signal bidirectional
flabel metal5 s 8920 848500 16920 856500 0 FreeSans 24000 0 0 0 vssio_5
port 124 nsew ground bidirectional
flabel metal5 s 8843 869500 16843 877500 0 FreeSans 24000 0 0 0 gpio5_3
port 125 nsew signal bidirectional
flabel metal5 s 8843 890500 16843 898500 0 FreeSans 24000 0 0 0 gpio5_2
port 126 nsew signal bidirectional
flabel metal5 s 8843 911500 16843 919500 0 FreeSans 24000 0 0 0 gpio5_1
port 127 nsew signal bidirectional
flabel metal5 s 8843 932500 16843 940500 0 FreeSans 24000 0 0 0 gpio5_0
port 128 nsew signal bidirectional
flabel metal5 s 8920 952500 16920 960500 0 FreeSans 24000 0 0 0 vssd2_1
port 129 nsew ground bidirectional
flabel metal5 s 8920 975500 16920 983500 0 FreeSans 24000 0 0 0 vddio_5
port 130 nsew power bidirectional
flabel metal3 s 47060 39793 51849 40793 0 FreeSans 8000 0 0 0 vccd0
port 131 nsew power bidirectional
flabel metal3 s 57100 39793 61902 40793 0 FreeSans 8000 0 0 0 vccd0
port 131 nsew power bidirectional
flabel metal3 s 206142 39793 210922 40793 0 FreeSans 8000 0 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 216121 39793 220901 40793 0 FreeSans 8000 0 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 228060 39793 232849 40793 0 FreeSans 8000 0 0 0 vssd0
port 133 nsew ground bidirectional
flabel metal3 s 238100 39793 242900 40793 0 FreeSans 8000 0 0 0 vssd0
port 133 nsew ground bidirectional
flabel metal3 s 338142 39793 342922 40793 0 FreeSans 8000 0 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 348121 39793 352901 40793 0 FreeSans 8000 0 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 364060 39793 368849 40793 0 FreeSans 8000 0 0 0 vccd0
port 131 nsew power bidirectional
flabel metal3 s 374100 39793 378902 40793 0 FreeSans 8000 0 0 0 vccd0
port 131 nsew power bidirectional
flabel metal3 s 478142 39793 482922 40793 0 FreeSans 8000 0 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 488121 39793 492901 40793 0 FreeSans 8000 0 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 500142 39793 504922 40793 0 FreeSans 8000 0 0 0 vssa3
port 135 nsew ground bidirectional
flabel metal3 s 510121 39793 514901 40793 0 FreeSans 8000 0 0 0 vssa3
port 135 nsew ground bidirectional
flabel metal3 s 526142 39793 530922 40793 0 FreeSans 8000 0 0 0 vdda3
port 136 nsew power bidirectional
flabel metal3 s 536121 39793 540901 40793 0 FreeSans 8000 0 0 0 vdda3
port 136 nsew power bidirectional
flabel metal3 s 552060 39793 556849 40793 0 FreeSans 8000 0 0 0 vssd0
port 133 nsew ground bidirectional
flabel metal3 s 562100 39793 566900 40793 0 FreeSans 8000 0 0 0 vssd0
port 133 nsew ground bidirectional
flabel metal3 s 676807 54742 677807 59522 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 676807 64721 677807 69501 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 676807 158660 677807 163449 0 FreeSans 8000 90 0 0 vssd1[0]
port 137 nsew ground bidirectional
flabel metal3 s 676807 168700 677807 173500 0 FreeSans 8000 90 0 0 vssd1[0]
port 137 nsew ground bidirectional
flabel metal3 s 676807 163749 677807 168400 0 FreeSans 8000 90 0 0 vccd1[0]
port 138 nsew power bidirectional
flabel metal3 s 676807 178742 677807 183522 0 FreeSans 8000 90 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 676807 188721 677807 193501 0 FreeSans 8000 90 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 676807 282742 677807 287522 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 676807 292721 677807 297501 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 676807 302742 677807 307522 0 FreeSans 8000 90 0 0 vdda1
port 139 nsew power bidirectional
flabel metal3 s 676807 312721 677807 317501 0 FreeSans 8000 90 0 0 vdda1
port 139 nsew power bidirectional
flabel metal3 s 676807 326742 677807 331522 0 FreeSans 8000 90 0 0 vssa1
port 140 nsew ground bidirectional
flabel metal3 s 676807 336721 677807 341501 0 FreeSans 8000 90 0 0 vssa1
port 140 nsew ground bidirectional
flabel metal3 s 676807 478660 677807 483449 0 FreeSans 8000 90 0 0 vccd1[1]
port 141 nsew power bidirectional
flabel metal3 s 676807 488700 677807 493502 0 FreeSans 8000 90 0 0 vccd1[1]
port 141 nsew power bidirectional
flabel metal3 s 676807 483748 677807 488410 0 FreeSans 8000 90 0 0 vssd1[1]
port 142 nsew ground bidirectional
flabel metal3 s 676807 523342 677807 528122 0 FreeSans 8000 90 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 676807 533321 677807 538101 0 FreeSans 8000 90 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 676807 675342 677807 680122 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 676807 685321 677807 690101 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 676807 695342 677807 700122 0 FreeSans 8000 90 0 0 vdda1
port 139 nsew power bidirectional
flabel metal3 s 676807 705321 677807 710101 0 FreeSans 8000 90 0 0 vdda1
port 139 nsew power bidirectional
flabel metal3 s 676807 719342 677807 724122 0 FreeSans 8000 90 0 0 vssa1
port 140 nsew ground bidirectional
flabel metal3 s 676807 729321 677807 734101 0 FreeSans 8000 90 0 0 vssa1
port 140 nsew ground bidirectional
flabel metal3 s 676807 739260 677807 744049 0 FreeSans 8000 90 0 0 vssd1[2]
port 143 nsew ground bidirectional
flabel metal3 s 676807 749300 677807 754100 0 FreeSans 8000 90 0 0 vssd1[2]
port 143 nsew ground bidirectional
flabel metal3 s 676807 744349 677807 749000 0 FreeSans 8000 90 0 0 vccd1[2]
port 144 nsew power bidirectional
flabel metal3 s 676807 843342 677807 848122 0 FreeSans 8000 90 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 676807 853321 677807 858101 0 FreeSans 8000 90 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 676807 947260 677807 952049 0 FreeSans 8000 90 0 0 vccd1[3]
port 145 nsew power bidirectional
flabel metal3 s 676807 957300 677807 962102 0 FreeSans 8000 90 0 0 vccd1[3]
port 145 nsew power bidirectional
flabel metal3 s 676807 952348 677807 957010 0 FreeSans 8000 90 0 0 vssd1[3]
port 146 nsew ground bidirectional
flabel metal3 s 676807 971342 677807 976122 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 676807 981321 677807 986101 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 668951 996807 673740 997807 0 FreeSans 8000 0 0 0 vssd1[4]
port 147 nsew ground bidirectional
flabel metal3 s 658900 996807 663700 997807 0 FreeSans 8000 0 0 0 vssd1[4]
port 147 nsew ground bidirectional
flabel metal3 s 664000 996807 668651 997807 0 FreeSans 8000 0 0 0 vccd1[4]
port 148 nsew power bidirectional
flabel metal3 s 549878 996807 554658 997807 0 FreeSans 8000 0 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 539899 996807 544679 997807 0 FreeSans 8000 0 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 526951 996807 531740 997807 0 FreeSans 8000 0 0 0 vccd1[5]
port 149 nsew power bidirectional
flabel metal3 s 516898 996807 521700 997807 0 FreeSans 8000 0 0 0 vccd1[5]
port 149 nsew power bidirectional
flabel metal3 s 521990 996807 526652 997807 0 FreeSans 8000 0 0 0 vssd1[5]
port 150 nsew ground bidirectional
flabel metal3 s 407878 996807 412658 997807 0 FreeSans 8000 0 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 397899 996807 402679 997807 0 FreeSans 8000 0 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 384878 996807 389658 997807 0 FreeSans 8000 0 0 0 vdda0
port 151 nsew power bidirectional
flabel metal3 s 374899 996807 379679 997807 0 FreeSans 8000 0 0 0 vdda0
port 151 nsew power bidirectional
flabel metal3 s 315878 996807 320658 997807 0 FreeSans 8000 0 0 0 vssa0
port 152 nsew ground bidirectional
flabel metal3 s 305899 996807 310679 997807 0 FreeSans 8000 0 0 0 vssa0
port 152 nsew ground bidirectional
flabel metal3 s 196951 996807 201740 997807 0 FreeSans 8000 0 0 0 vssd2[0]
port 153 nsew ground bidirectional
flabel metal3 s 186900 996807 191700 997807 0 FreeSans 8000 0 0 0 vssd2[0]
port 153 nsew ground bidirectional
flabel metal3 s 192000 996807 196651 997807 0 FreeSans 8000 0 0 0 vccd2[0]
port 154 nsew power bidirectional
flabel metal3 s 173878 996807 178658 997807 0 FreeSans 8000 0 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 163899 996807 168679 997807 0 FreeSans 8000 0 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 54951 996807 59740 997807 0 FreeSans 8000 0 0 0 vccd2[1]
port 155 nsew power bidirectional
flabel metal3 s 44898 996807 49700 997807 0 FreeSans 8000 0 0 0 vccd2[1]
port 155 nsew power bidirectional
flabel metal3 s 49990 996807 54652 997807 0 FreeSans 8000 0 0 0 vssd2[1]
port 156 nsew ground bidirectional
flabel metal3 s 39793 972099 40793 976879 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 39793 982078 40793 986858 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 39793 949100 40793 953900 0 FreeSans 8000 90 0 0 vssd2[2]
port 157 nsew ground bidirectional
flabel metal3 s 39793 959151 40793 963940 0 FreeSans 8000 90 0 0 vssd2[2]
port 157 nsew ground bidirectional
flabel metal3 s 39793 845099 40793 849879 0 FreeSans 8000 90 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 39793 855078 40793 859858 0 FreeSans 8000 90 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 39793 741098 40793 745900 0 FreeSans 8000 90 0 0 vccd2[3]
port 159 nsew power bidirectional
flabel metal3 s 39793 751151 40793 755940 0 FreeSans 8000 90 0 0 vccd2[3]
port 159 nsew power bidirectional
flabel metal3 s 39793 746190 40793 750852 0 FreeSans 8000 90 0 0 vssd2[3]
port 160 nsew ground bidirectional
flabel metal3 s 39793 721099 40793 725879 0 FreeSans 8000 90 0 0 vssa2
port 161 nsew ground bidirectional
flabel metal3 s 39793 731078 40793 735858 0 FreeSans 8000 90 0 0 vssa2
port 161 nsew ground bidirectional
flabel metal3 s 39793 698099 40793 702879 0 FreeSans 8000 90 0 0 vdda2
port 162 nsew power bidirectional
flabel metal3 s 39793 708078 40793 712858 0 FreeSans 8000 90 0 0 vdda2
port 162 nsew power bidirectional
flabel metal3 s 39793 678099 40793 682879 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 39793 688078 40793 692858 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 39793 526099 40793 530879 0 FreeSans 8000 90 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 39793 536078 40793 540858 0 FreeSans 8000 90 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 39793 481500 40793 486300 0 FreeSans 8000 90 0 0 vssd2[4]
port 163 nsew ground bidirectional
flabel metal3 s 39793 491551 40793 496340 0 FreeSans 8000 90 0 0 vssd2[4]
port 163 nsew ground bidirectional
flabel metal3 s 39793 486600 40793 491251 0 FreeSans 8000 90 0 0 vccd2[4]
port 164 nsew power bidirectional
flabel metal3 s 39793 329499 40793 334279 0 FreeSans 8000 90 0 0 vssa2
port 161 nsew ground bidirectional
flabel metal3 s 39793 339478 40793 344258 0 FreeSans 8000 90 0 0 vssa2
port 161 nsew ground bidirectional
flabel metal3 s 39793 306499 40793 311279 0 FreeSans 8000 90 0 0 vdda2
port 162 nsew power bidirectional
flabel metal3 s 39793 316478 40793 321258 0 FreeSans 8000 90 0 0 vdda2
port 162 nsew power bidirectional
flabel metal3 s 39793 286499 40793 291279 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 39793 296478 40793 301258 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 39793 182499 40793 187279 0 FreeSans 8000 90 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 39793 192478 40793 197258 0 FreeSans 8000 90 0 0 vssio
port 132 nsew ground bidirectional
flabel metal3 s 39793 159498 40793 164300 0 FreeSans 8000 90 0 0 vccd2[5]
port 165 nsew power bidirectional
flabel metal3 s 39793 169551 40793 174340 0 FreeSans 8000 90 0 0 vccd2[5]
port 165 nsew power bidirectional
flabel metal3 s 39793 164590 40793 169252 0 FreeSans 8000 90 0 0 vssd2[5]
port 166 nsew ground bidirectional
flabel metal3 s 39793 55499 40793 60279 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal3 s 39793 65478 40793 70258 0 FreeSans 8000 90 0 0 vddio
port 134 nsew power bidirectional
flabel metal2 s 68457 40710 68509 40910 0 FreeSans 320 90 0 0 select_tie_lo_esd
port 167 nsew signal output
flabel metal2 s 68757 40710 68809 40910 0 FreeSans 320 90 0 0 select_in
port 168 nsew signal output
flabel metal2 s 69059 40710 69111 40910 0 FreeSans 320 90 0 0 select_tie_hi_esd
port 169 nsew signal output
flabel metal2 s 69357 40710 69409 40910 0 FreeSans 320 90 0 0 select_enable_vddio
port 170 nsew signal input
flabel metal2 s 69657 40710 69709 40910 0 FreeSans 320 90 0 0 select_slow
port 171 nsew signal input
flabel metal2 s 69957 40710 70085 40910 0 FreeSans 320 90 0 0 select_pad_a_esd_0_h
port 172 nsew signal bidirectional
flabel metal2 s 71215 40710 71345 40910 0 FreeSans 320 90 0 0 select_pad_a_esd_1_h
port 173 nsew signal bidirectional
flabel metal2 s 72223 40710 72437 40910 0 FreeSans 320 90 0 0 select_pad_a_noesd_h
port 174 nsew signal bidirectional
flabel metal2 s 72689 40710 72741 40910 0 FreeSans 320 90 0 0 select_analog_en
port 175 nsew signal input
flabel metal2 s 75603 40710 75655 40910 0 FreeSans 320 90 0 0 select_analog_pol
port 176 nsew signal input
flabel metal2 s 75899 40710 75951 40910 0 FreeSans 320 90 0 0 select_inp_dis
port 177 nsew signal input
flabel metal2 s 77270 40710 77326 40910 0 FreeSans 320 90 0 0 select_enable_inp_h
port 178 nsew signal input
flabel metal2 s 77856 40710 77908 40910 0 FreeSans 320 90 0 0 select_enable_h
port 179 nsew signal input
flabel metal2 s 78585 40710 78637 40910 0 FreeSans 320 90 0 0 select_hld_h_n
port 180 nsew signal input
flabel metal2 s 78899 40710 78951 40910 0 FreeSans 320 90 0 0 select_analog_sel
port 181 nsew signal input
flabel metal2 s 79250 40710 79302 40910 0 FreeSans 320 90 0 0 select_dm[2]
port 182 nsew signal input
flabel metal2 s 71581 40710 71633 40910 0 FreeSans 320 90 0 0 select_dm[1]
port 183 nsew signal input
flabel metal2 s 74977 40710 75029 40910 0 FreeSans 320 90 0 0 select_dm[0]
port 184 nsew signal input
flabel metal2 s 79628 40710 79680 40910 0 FreeSans 320 90 0 0 select_hld_ovr
port 185 nsew signal input
flabel metal2 s 80477 40710 80529 40910 0 FreeSans 320 90 0 0 select_out
port 186 nsew signal input
flabel metal2 s 81686 40710 81738 40910 0 FreeSans 320 90 0 0 select_enable_vswitch_h
port 187 nsew signal input
flabel metal2 s 82397 40710 82449 40910 0 FreeSans 320 90 0 0 select_enable_vdda_h
port 188 nsew signal input
flabel metal2 s 83645 40710 83697 40910 0 FreeSans 320 90 0 0 select_vtrip_sel
port 189 nsew signal input
flabel metal2 s 83965 40710 84017 40910 0 FreeSans 320 90 0 0 select_ib_mode_sel
port 190 nsew signal input
flabel metal2 s 84279 40710 84331 40910 0 FreeSans 320 90 0 0 select_oe_n
port 191 nsew signal input
flabel metal2 s 84797 40710 84921 40910 0 FreeSans 320 90 0 0 select_in_h
port 192 nsew signal input
flabel metal2 s 67493 40710 67545 40910 0 FreeSans 320 90 0 0 select_zero
port 193 nsew signal output
flabel metal2 s 67131 40710 67183 40910 0 FreeSans 320 90 0 0 select_one
port 194 nsew signal output
flabel metal2 s 92353 40300 92557 40600 0 FreeSans 320 90 0 0 resetb_tie_weak_hi_h
port 195 nsew signal output
flabel metal2 s 100396 40300 100448 40600 0 FreeSans 320 90 0 0 resetb_disable_pullup_h
port 196 nsew signal input
flabel metal2 s 100769 40300 100899 40600 0 FreeSans 320 90 0 0 resetb_tie_hi_esd
port 197 nsew signal output
flabel metal2 s 101067 40300 101213 40600 0 FreeSans 320 90 0 0 resetb_xres_h_n
port 198 nsew signal output
flabel metal2 s 101354 40300 101484 40600 0 FreeSans 320 90 0 0 resetb_tie_lo_esd
port 199 nsew signal output
flabel metal2 s 101969 40330 102023 40600 0 FreeSans 320 90 0 0 resetb_inp_sel_h
port 200 nsew signal input
flabel metal2 s 102468 40300 102528 40600 0 FreeSans 320 90 0 0 resetb_en_vddio_sig_h
port 201 nsew signal input
flabel metal2 s 102755 40300 102985 40600 0 FreeSans 320 90 0 0 resetb_filt_in_h
port 202 nsew signal input
flabel metal2 s 103218 40300 103551 40600 0 FreeSans 320 90 0 0 resetb_pad_a_esd_h
port 203 nsew signal output
flabel metal2 s 103973 40300 104089 40600 0 FreeSans 320 90 0 0 resetb_pullup_h
port 204 nsew signal input
flabel metal2 s 104491 40300 104543 40600 0 FreeSans 320 90 0 0 resetb_enable_h
port 205 nsew signal input
flabel metal2 s 105221 40300 105315 40600 0 FreeSans 320 90 0 0 resetb_enable_vddio
port 206 nsew signal input
flabel metal2 s 113457 40710 113509 40910 0 FreeSans 320 90 0 0 gpio8_0_tie_lo_esd
port 207 nsew signal output
flabel metal2 s 113757 40710 113809 40910 0 FreeSans 320 90 0 0 gpio8_0_in
port 208 nsew signal output
flabel metal2 s 114059 40710 114111 40910 0 FreeSans 320 90 0 0 gpio8_0_tie_hi_esd
port 209 nsew signal output
flabel metal2 s 114357 40710 114409 40910 0 FreeSans 320 90 0 0 gpio8_0_enable_vddio
port 210 nsew signal input
flabel metal2 s 114657 40710 114709 40910 0 FreeSans 320 90 0 0 gpio8_0_slow
port 211 nsew signal input
flabel metal2 s 114957 40710 115085 40910 0 FreeSans 320 90 0 0 gpio8_0_pad_a_esd_0_h
port 212 nsew signal bidirectional
flabel metal2 s 116215 40710 116345 40910 0 FreeSans 320 90 0 0 gpio8_0_pad_a_esd_1_h
port 213 nsew signal bidirectional
flabel metal2 s 117223 40710 117437 40910 0 FreeSans 320 90 0 0 gpio8_0_pad_a_noesd_h
port 214 nsew signal bidirectional
flabel metal2 s 117689 40710 117741 40910 0 FreeSans 320 90 0 0 gpio8_0_analog_en
port 215 nsew signal input
flabel metal2 s 120603 40710 120655 40910 0 FreeSans 320 90 0 0 gpio8_0_analog_pol
port 216 nsew signal input
flabel metal2 s 120899 40710 120951 40910 0 FreeSans 320 90 0 0 gpio8_0_inp_dis
port 217 nsew signal input
flabel metal2 s 122270 40710 122326 40910 0 FreeSans 320 90 0 0 gpio8_0_enable_inp_h
port 218 nsew signal input
flabel metal2 s 122856 40710 122908 40910 0 FreeSans 320 90 0 0 gpio8_0_enable_h
port 219 nsew signal input
flabel metal2 s 123585 40710 123637 40910 0 FreeSans 320 90 0 0 gpio8_0_hld_h_n
port 220 nsew signal input
flabel metal2 s 123899 40710 123951 40910 0 FreeSans 320 90 0 0 gpio8_0_analog_sel
port 221 nsew signal input
flabel metal2 s 124250 40710 124302 40910 0 FreeSans 320 90 0 0 gpio8_0_dm[2]
port 222 nsew signal input
flabel metal2 s 116581 40710 116633 40910 0 FreeSans 320 90 0 0 gpio8_0_dm[1]
port 223 nsew signal input
flabel metal2 s 119977 40710 120029 40910 0 FreeSans 320 90 0 0 gpio8_0_dm[0]
port 224 nsew signal input
flabel metal2 s 124628 40710 124680 40910 0 FreeSans 320 90 0 0 gpio8_0_hld_ovr
port 225 nsew signal input
flabel metal2 s 125477 40710 125529 40910 0 FreeSans 320 90 0 0 gpio8_0_out
port 226 nsew signal input
flabel metal2 s 126686 40710 126738 40910 0 FreeSans 320 90 0 0 gpio8_0_enable_vswitch_h
port 227 nsew signal input
flabel metal2 s 127397 40710 127449 40910 0 FreeSans 320 90 0 0 gpio8_0_enable_vdda_h
port 228 nsew signal input
flabel metal2 s 128645 40710 128697 40910 0 FreeSans 320 90 0 0 gpio8_0_vtrip_sel
port 229 nsew signal input
flabel metal2 s 128965 40710 129017 40910 0 FreeSans 320 90 0 0 gpio8_0_ib_mode_sel
port 230 nsew signal input
flabel metal2 s 129279 40710 129331 40910 0 FreeSans 320 90 0 0 gpio8_0_oe_n
port 231 nsew signal input
flabel metal2 s 129797 40710 129921 40910 0 FreeSans 320 90 0 0 gpio8_0_in_h
port 232 nsew signal input
flabel metal2 s 112493 40710 112545 40910 0 FreeSans 320 90 0 0 gpio8_0_zero
port 233 nsew signal output
flabel metal2 s 112131 40710 112183 40910 0 FreeSans 320 90 0 0 gpio8_0_one
port 234 nsew signal output
flabel metal2 s 136457 40710 136509 40910 0 FreeSans 320 90 0 0 gpio8_1_tie_lo_esd
port 235 nsew signal output
flabel metal2 s 136757 40710 136809 40910 0 FreeSans 320 90 0 0 gpio8_1_in
port 236 nsew signal output
flabel metal2 s 137059 40710 137111 40910 0 FreeSans 320 90 0 0 gpio8_1_tie_hi_esd
port 237 nsew signal output
flabel metal2 s 137357 40710 137409 40910 0 FreeSans 320 90 0 0 gpio8_1_enable_vddio
port 238 nsew signal input
flabel metal2 s 137657 40710 137709 40910 0 FreeSans 320 90 0 0 gpio8_1_slow
port 239 nsew signal input
flabel metal2 s 137957 40710 138085 40910 0 FreeSans 320 90 0 0 gpio8_1_pad_a_esd_0_h
port 240 nsew signal bidirectional
flabel metal2 s 139215 40710 139345 40910 0 FreeSans 320 90 0 0 gpio8_1_pad_a_esd_1_h
port 241 nsew signal bidirectional
flabel metal2 s 140223 40710 140437 40910 0 FreeSans 320 90 0 0 gpio8_1_pad_a_noesd_h
port 242 nsew signal bidirectional
flabel metal2 s 140689 40710 140741 40910 0 FreeSans 320 90 0 0 gpio8_1_analog_en
port 243 nsew signal input
flabel metal2 s 143603 40710 143655 40910 0 FreeSans 320 90 0 0 gpio8_1_analog_pol
port 244 nsew signal input
flabel metal2 s 143899 40710 143951 40910 0 FreeSans 320 90 0 0 gpio8_1_inp_dis
port 245 nsew signal input
flabel metal2 s 145270 40710 145326 40910 0 FreeSans 320 90 0 0 gpio8_1_enable_inp_h
port 246 nsew signal input
flabel metal2 s 145856 40710 145908 40910 0 FreeSans 320 90 0 0 gpio8_1_enable_h
port 247 nsew signal input
flabel metal2 s 146585 40710 146637 40910 0 FreeSans 320 90 0 0 gpio8_1_hld_h_n
port 248 nsew signal input
flabel metal2 s 146899 40710 146951 40910 0 FreeSans 320 90 0 0 gpio8_1_analog_sel
port 249 nsew signal input
flabel metal2 s 147250 40710 147302 40910 0 FreeSans 320 90 0 0 gpio8_1_dm[2]
port 250 nsew signal input
flabel metal2 s 139581 40710 139633 40910 0 FreeSans 320 90 0 0 gpio8_1_dm[1]
port 251 nsew signal input
flabel metal2 s 142977 40710 143029 40910 0 FreeSans 320 90 0 0 gpio8_1_dm[0]
port 252 nsew signal input
flabel metal2 s 147628 40710 147680 40910 0 FreeSans 320 90 0 0 gpio8_1_hld_ovr
port 253 nsew signal input
flabel metal2 s 148477 40710 148529 40910 0 FreeSans 320 90 0 0 gpio8_1_out
port 254 nsew signal input
flabel metal2 s 149686 40710 149738 40910 0 FreeSans 320 90 0 0 gpio8_1_enable_vswitch_h
port 255 nsew signal input
flabel metal2 s 150397 40710 150449 40910 0 FreeSans 320 90 0 0 gpio8_1_enable_vdda_h
port 256 nsew signal input
flabel metal2 s 151645 40710 151697 40910 0 FreeSans 320 90 0 0 gpio8_1_vtrip_sel
port 257 nsew signal input
flabel metal2 s 151965 40710 152017 40910 0 FreeSans 320 90 0 0 gpio8_1_ib_mode_sel
port 258 nsew signal input
flabel metal2 s 152279 40710 152331 40910 0 FreeSans 320 90 0 0 gpio8_1_oe_n
port 259 nsew signal input
flabel metal2 s 152797 40710 152921 40910 0 FreeSans 320 90 0 0 gpio8_1_in_h
port 260 nsew signal input
flabel metal2 s 135493 40710 135545 40910 0 FreeSans 320 90 0 0 gpio8_1_zero
port 261 nsew signal output
flabel metal2 s 135131 40710 135183 40910 0 FreeSans 320 90 0 0 gpio8_1_one
port 262 nsew signal output
flabel metal2 s 159457 40710 159509 40910 0 FreeSans 320 90 0 0 gpio8_2_tie_lo_esd
port 263 nsew signal output
flabel metal2 s 159757 40710 159809 40910 0 FreeSans 320 90 0 0 gpio8_2_in
port 264 nsew signal output
flabel metal2 s 160059 40710 160111 40910 0 FreeSans 320 90 0 0 gpio8_2_tie_hi_esd
port 265 nsew signal output
flabel metal2 s 160357 40710 160409 40910 0 FreeSans 320 90 0 0 gpio8_2_enable_vddio
port 266 nsew signal input
flabel metal2 s 160657 40710 160709 40910 0 FreeSans 320 90 0 0 gpio8_2_slow
port 267 nsew signal input
flabel metal2 s 160957 40710 161085 40910 0 FreeSans 320 90 0 0 gpio8_2_pad_a_esd_0_h
port 268 nsew signal bidirectional
flabel metal2 s 162215 40710 162345 40910 0 FreeSans 320 90 0 0 gpio8_2_pad_a_esd_1_h
port 269 nsew signal bidirectional
flabel metal2 s 163223 40710 163437 40910 0 FreeSans 320 90 0 0 gpio8_2_pad_a_noesd_h
port 270 nsew signal bidirectional
flabel metal2 s 163689 40710 163741 40910 0 FreeSans 320 90 0 0 gpio8_2_analog_en
port 271 nsew signal input
flabel metal2 s 166603 40710 166655 40910 0 FreeSans 320 90 0 0 gpio8_2_analog_pol
port 272 nsew signal input
flabel metal2 s 166899 40710 166951 40910 0 FreeSans 320 90 0 0 gpio8_2_inp_dis
port 273 nsew signal input
flabel metal2 s 168270 40710 168326 40910 0 FreeSans 320 90 0 0 gpio8_2_enable_inp_h
port 274 nsew signal input
flabel metal2 s 168856 40710 168908 40910 0 FreeSans 320 90 0 0 gpio8_2_enable_h
port 275 nsew signal input
flabel metal2 s 169585 40710 169637 40910 0 FreeSans 320 90 0 0 gpio8_2_hld_h_n
port 276 nsew signal input
flabel metal2 s 169899 40710 169951 40910 0 FreeSans 320 90 0 0 gpio8_2_analog_sel
port 277 nsew signal input
flabel metal2 s 170250 40710 170302 40910 0 FreeSans 320 90 0 0 gpio8_2_dm[2]
port 278 nsew signal input
flabel metal2 s 162581 40710 162633 40910 0 FreeSans 320 90 0 0 gpio8_2_dm[1]
port 279 nsew signal input
flabel metal2 s 165977 40710 166029 40910 0 FreeSans 320 90 0 0 gpio8_2_dm[0]
port 280 nsew signal input
flabel metal2 s 170628 40710 170680 40910 0 FreeSans 320 90 0 0 gpio8_2_hld_ovr
port 281 nsew signal input
flabel metal2 s 171477 40710 171529 40910 0 FreeSans 320 90 0 0 gpio8_2_out
port 282 nsew signal input
flabel metal2 s 172686 40710 172738 40910 0 FreeSans 320 90 0 0 gpio8_2_enable_vswitch_h
port 283 nsew signal input
flabel metal2 s 173397 40710 173449 40910 0 FreeSans 320 90 0 0 gpio8_2_enable_vdda_h
port 284 nsew signal input
flabel metal2 s 174645 40710 174697 40910 0 FreeSans 320 90 0 0 gpio8_2_vtrip_sel
port 285 nsew signal input
flabel metal2 s 174965 40710 175017 40910 0 FreeSans 320 90 0 0 gpio8_2_ib_mode_sel
port 286 nsew signal input
flabel metal2 s 175279 40710 175331 40910 0 FreeSans 320 90 0 0 gpio8_2_oe_n
port 287 nsew signal input
flabel metal2 s 175797 40710 175921 40910 0 FreeSans 320 90 0 0 gpio8_2_in_h
port 288 nsew signal input
flabel metal2 s 158493 40710 158545 40910 0 FreeSans 320 90 0 0 gpio8_2_zero
port 289 nsew signal output
flabel metal2 s 158131 40710 158183 40910 0 FreeSans 320 90 0 0 gpio8_2_one
port 290 nsew signal output
flabel metal2 s 182457 40710 182509 40910 0 FreeSans 320 90 0 0 gpio8_3_tie_lo_esd
port 291 nsew signal output
flabel metal2 s 182757 40710 182809 40910 0 FreeSans 320 90 0 0 gpio8_3_in
port 292 nsew signal output
flabel metal2 s 183059 40710 183111 40910 0 FreeSans 320 90 0 0 gpio8_3_tie_hi_esd
port 293 nsew signal output
flabel metal2 s 183357 40710 183409 40910 0 FreeSans 320 90 0 0 gpio8_3_enable_vddio
port 294 nsew signal input
flabel metal2 s 183657 40710 183709 40910 0 FreeSans 320 90 0 0 gpio8_3_slow
port 295 nsew signal input
flabel metal2 s 183957 40710 184085 40910 0 FreeSans 320 90 0 0 gpio8_3_pad_a_esd_0_h
port 296 nsew signal bidirectional
flabel metal2 s 185215 40710 185345 40910 0 FreeSans 320 90 0 0 gpio8_3_pad_a_esd_1_h
port 297 nsew signal bidirectional
flabel metal2 s 186223 40710 186437 40910 0 FreeSans 320 90 0 0 gpio8_3_pad_a_noesd_h
port 298 nsew signal bidirectional
flabel metal2 s 186689 40710 186741 40910 0 FreeSans 320 90 0 0 gpio8_3_analog_en
port 299 nsew signal input
flabel metal2 s 189603 40710 189655 40910 0 FreeSans 320 90 0 0 gpio8_3_analog_pol
port 300 nsew signal input
flabel metal2 s 189899 40710 189951 40910 0 FreeSans 320 90 0 0 gpio8_3_inp_dis
port 301 nsew signal input
flabel metal2 s 191270 40710 191326 40910 0 FreeSans 320 90 0 0 gpio8_3_enable_inp_h
port 302 nsew signal input
flabel metal2 s 191856 40710 191908 40910 0 FreeSans 320 90 0 0 gpio8_3_enable_h
port 303 nsew signal input
flabel metal2 s 192585 40710 192637 40910 0 FreeSans 320 90 0 0 gpio8_3_hld_h_n
port 304 nsew signal input
flabel metal2 s 192899 40710 192951 40910 0 FreeSans 320 90 0 0 gpio8_3_analog_sel
port 305 nsew signal input
flabel metal2 s 193250 40710 193302 40910 0 FreeSans 320 90 0 0 gpio8_3_dm[2]
port 306 nsew signal input
flabel metal2 s 185581 40710 185633 40910 0 FreeSans 320 90 0 0 gpio8_3_dm[1]
port 307 nsew signal input
flabel metal2 s 188977 40710 189029 40910 0 FreeSans 320 90 0 0 gpio8_3_dm[0]
port 308 nsew signal input
flabel metal2 s 193628 40710 193680 40910 0 FreeSans 320 90 0 0 gpio8_3_hld_ovr
port 309 nsew signal input
flabel metal2 s 194477 40710 194529 40910 0 FreeSans 320 90 0 0 gpio8_3_out
port 310 nsew signal input
flabel metal2 s 195686 40710 195738 40910 0 FreeSans 320 90 0 0 gpio8_3_enable_vswitch_h
port 311 nsew signal input
flabel metal2 s 196397 40710 196449 40910 0 FreeSans 320 90 0 0 gpio8_3_enable_vdda_h
port 312 nsew signal input
flabel metal2 s 197645 40710 197697 40910 0 FreeSans 320 90 0 0 gpio8_3_vtrip_sel
port 313 nsew signal input
flabel metal2 s 197965 40710 198017 40910 0 FreeSans 320 90 0 0 gpio8_3_ib_mode_sel
port 314 nsew signal input
flabel metal2 s 198279 40710 198331 40910 0 FreeSans 320 90 0 0 gpio8_3_oe_n
port 315 nsew signal input
flabel metal2 s 198797 40710 198921 40910 0 FreeSans 320 90 0 0 gpio8_3_in_h
port 316 nsew signal input
flabel metal2 s 181493 40710 181545 40910 0 FreeSans 320 90 0 0 gpio8_3_zero
port 317 nsew signal output
flabel metal2 s 181131 40710 181183 40910 0 FreeSans 320 90 0 0 gpio8_3_one
port 318 nsew signal output
flabel metal2 s 255438 40600 257234 41000 0 FreeSans 320 0 0 0 xi0_core
port 319 nsew analog bidirectional
flabel metal2 s 277438 40600 279234 41000 0 FreeSans 320 0 0 0 xo0_core
port 320 nsew analog bidirectional
flabel metal2 s 299438 40600 301234 41000 0 FreeSans 320 0 0 0 xi1_core
port 321 nsew analog bidirectional
flabel metal2 s 321438 40600 323234 41000 0 FreeSans 320 0 0 0 xo1_core
port 322 nsew analog bidirectional
flabel metal2 s 385457 40710 385509 40910 0 FreeSans 320 90 0 0 gpio8_4_tie_lo_esd
port 323 nsew signal output
flabel metal2 s 385757 40710 385809 40910 0 FreeSans 320 90 0 0 gpio8_4_in
port 324 nsew signal output
flabel metal2 s 386059 40710 386111 40910 0 FreeSans 320 90 0 0 gpio8_4_tie_hi_esd
port 325 nsew signal output
flabel metal2 s 386357 40710 386409 40910 0 FreeSans 320 90 0 0 gpio8_4_enable_vddio
port 326 nsew signal input
flabel metal2 s 386657 40710 386709 40910 0 FreeSans 320 90 0 0 gpio8_4_slow
port 327 nsew signal input
flabel metal2 s 386957 40710 387085 40910 0 FreeSans 320 90 0 0 gpio8_4_pad_a_esd_0_h
port 328 nsew signal bidirectional
flabel metal2 s 388215 40710 388345 40910 0 FreeSans 320 90 0 0 gpio8_4_pad_a_esd_1_h
port 329 nsew signal bidirectional
flabel metal2 s 389223 40710 389437 40910 0 FreeSans 320 90 0 0 gpio8_4_pad_a_noesd_h
port 330 nsew signal bidirectional
flabel metal2 s 389689 40710 389741 40910 0 FreeSans 320 90 0 0 gpio8_4_analog_en
port 331 nsew signal input
flabel metal2 s 392603 40710 392655 40910 0 FreeSans 320 90 0 0 gpio8_4_analog_pol
port 332 nsew signal input
flabel metal2 s 392899 40710 392951 40910 0 FreeSans 320 90 0 0 gpio8_4_inp_dis
port 333 nsew signal input
flabel metal2 s 394270 40710 394326 40910 0 FreeSans 320 90 0 0 gpio8_4_enable_inp_h
port 334 nsew signal input
flabel metal2 s 394856 40710 394908 40910 0 FreeSans 320 90 0 0 gpio8_4_enable_h
port 335 nsew signal input
flabel metal2 s 395585 40710 395637 40910 0 FreeSans 320 90 0 0 gpio8_4_hld_h_n
port 336 nsew signal input
flabel metal2 s 395899 40710 395951 40910 0 FreeSans 320 90 0 0 gpio8_4_analog_sel
port 337 nsew signal input
flabel metal2 s 396250 40710 396302 40910 0 FreeSans 320 90 0 0 gpio8_4_dm[2]
port 338 nsew signal input
flabel metal2 s 388581 40710 388633 40910 0 FreeSans 320 90 0 0 gpio8_4_dm[1]
port 339 nsew signal input
flabel metal2 s 391977 40710 392029 40910 0 FreeSans 320 90 0 0 gpio8_4_dm[0]
port 340 nsew signal input
flabel metal2 s 396628 40710 396680 40910 0 FreeSans 320 90 0 0 gpio8_4_hld_ovr
port 341 nsew signal input
flabel metal2 s 397477 40710 397529 40910 0 FreeSans 320 90 0 0 gpio8_4_out
port 342 nsew signal input
flabel metal2 s 398686 40710 398738 40910 0 FreeSans 320 90 0 0 gpio8_4_enable_vswitch_h
port 343 nsew signal input
flabel metal2 s 399397 40710 399449 40910 0 FreeSans 320 90 0 0 gpio8_4_enable_vdda_h
port 344 nsew signal input
flabel metal2 s 400645 40710 400697 40910 0 FreeSans 320 90 0 0 gpio8_4_vtrip_sel
port 345 nsew signal input
flabel metal2 s 400965 40710 401017 40910 0 FreeSans 320 90 0 0 gpio8_4_ib_mode_sel
port 346 nsew signal input
flabel metal2 s 401279 40710 401331 40910 0 FreeSans 320 90 0 0 gpio8_4_oe_n
port 347 nsew signal input
flabel metal2 s 401797 40710 401921 40910 0 FreeSans 320 90 0 0 gpio8_4_in_h
port 348 nsew signal input
flabel metal2 s 384493 40710 384545 40910 0 FreeSans 320 90 0 0 gpio8_4_zero
port 349 nsew signal output
flabel metal2 s 384131 40710 384183 40910 0 FreeSans 320 90 0 0 gpio8_4_one
port 350 nsew signal output
flabel metal2 s 408457 40710 408509 40910 0 FreeSans 320 90 0 0 gpio8_5_tie_lo_esd
port 351 nsew signal output
flabel metal2 s 408757 40710 408809 40910 0 FreeSans 320 90 0 0 gpio8_5_in
port 352 nsew signal output
flabel metal2 s 409059 40710 409111 40910 0 FreeSans 320 90 0 0 gpio8_5_tie_hi_esd
port 353 nsew signal output
flabel metal2 s 409357 40710 409409 40910 0 FreeSans 320 90 0 0 gpio8_5_enable_vddio
port 354 nsew signal input
flabel metal2 s 409657 40710 409709 40910 0 FreeSans 320 90 0 0 gpio8_5_slow
port 355 nsew signal input
flabel metal2 s 409957 40710 410085 40910 0 FreeSans 320 90 0 0 gpio8_5_pad_a_esd_0_h
port 356 nsew signal bidirectional
flabel metal2 s 411215 40710 411345 40910 0 FreeSans 320 90 0 0 gpio8_5_pad_a_esd_1_h
port 357 nsew signal bidirectional
flabel metal2 s 412223 40710 412437 40910 0 FreeSans 320 90 0 0 gpio8_5_pad_a_noesd_h
port 358 nsew signal bidirectional
flabel metal2 s 412689 40710 412741 40910 0 FreeSans 320 90 0 0 gpio8_5_analog_en
port 359 nsew signal input
flabel metal2 s 415603 40710 415655 40910 0 FreeSans 320 90 0 0 gpio8_5_analog_pol
port 360 nsew signal input
flabel metal2 s 415899 40710 415951 40910 0 FreeSans 320 90 0 0 gpio8_5_inp_dis
port 361 nsew signal input
flabel metal2 s 417270 40710 417326 40910 0 FreeSans 320 90 0 0 gpio8_5_enable_inp_h
port 362 nsew signal input
flabel metal2 s 417856 40710 417908 40910 0 FreeSans 320 90 0 0 gpio8_5_enable_h
port 363 nsew signal input
flabel metal2 s 418585 40710 418637 40910 0 FreeSans 320 90 0 0 gpio8_5_hld_h_n
port 364 nsew signal input
flabel metal2 s 418899 40710 418951 40910 0 FreeSans 320 90 0 0 gpio8_5_analog_sel
port 365 nsew signal input
flabel metal2 s 419250 40710 419302 40910 0 FreeSans 320 90 0 0 gpio8_5_dm[2]
port 366 nsew signal input
flabel metal2 s 411581 40710 411633 40910 0 FreeSans 320 90 0 0 gpio8_5_dm[1]
port 367 nsew signal input
flabel metal2 s 414977 40710 415029 40910 0 FreeSans 320 90 0 0 gpio8_5_dm[0]
port 368 nsew signal input
flabel metal2 s 419628 40710 419680 40910 0 FreeSans 320 90 0 0 gpio8_5_hld_ovr
port 369 nsew signal input
flabel metal2 s 420477 40710 420529 40910 0 FreeSans 320 90 0 0 gpio8_5_out
port 370 nsew signal input
flabel metal2 s 421686 40710 421738 40910 0 FreeSans 320 90 0 0 gpio8_5_enable_vswitch_h
port 371 nsew signal input
flabel metal2 s 422397 40710 422449 40910 0 FreeSans 320 90 0 0 gpio8_5_enable_vdda_h
port 372 nsew signal input
flabel metal2 s 423645 40710 423697 40910 0 FreeSans 320 90 0 0 gpio8_5_vtrip_sel
port 373 nsew signal input
flabel metal2 s 423965 40710 424017 40910 0 FreeSans 320 90 0 0 gpio8_5_ib_mode_sel
port 374 nsew signal input
flabel metal2 s 424279 40710 424331 40910 0 FreeSans 320 90 0 0 gpio8_5_oe_n
port 375 nsew signal input
flabel metal2 s 424797 40710 424921 40910 0 FreeSans 320 90 0 0 gpio8_5_in_h
port 376 nsew signal input
flabel metal2 s 407493 40710 407545 40910 0 FreeSans 320 90 0 0 gpio8_5_zero
port 377 nsew signal output
flabel metal2 s 407131 40710 407183 40910 0 FreeSans 320 90 0 0 gpio8_5_one
port 378 nsew signal output
flabel metal2 s 431457 40710 431509 40910 0 FreeSans 320 90 0 0 gpio8_6_tie_lo_esd
port 379 nsew signal output
flabel metal2 s 431757 40710 431809 40910 0 FreeSans 320 90 0 0 gpio8_6_in
port 380 nsew signal output
flabel metal2 s 432059 40710 432111 40910 0 FreeSans 320 90 0 0 gpio8_6_tie_hi_esd
port 381 nsew signal output
flabel metal2 s 432357 40710 432409 40910 0 FreeSans 320 90 0 0 gpio8_6_enable_vddio
port 382 nsew signal input
flabel metal2 s 432657 40710 432709 40910 0 FreeSans 320 90 0 0 gpio8_6_slow
port 383 nsew signal input
flabel metal2 s 432957 40710 433085 40910 0 FreeSans 320 90 0 0 gpio8_6_pad_a_esd_0_h
port 384 nsew signal bidirectional
flabel metal2 s 434215 40710 434345 40910 0 FreeSans 320 90 0 0 gpio8_6_pad_a_esd_1_h
port 385 nsew signal bidirectional
flabel metal2 s 435223 40710 435437 40910 0 FreeSans 320 90 0 0 gpio8_6_pad_a_noesd_h
port 386 nsew signal bidirectional
flabel metal2 s 435689 40710 435741 40910 0 FreeSans 320 90 0 0 gpio8_6_analog_en
port 387 nsew signal input
flabel metal2 s 438603 40710 438655 40910 0 FreeSans 320 90 0 0 gpio8_6_analog_pol
port 388 nsew signal input
flabel metal2 s 438899 40710 438951 40910 0 FreeSans 320 90 0 0 gpio8_6_inp_dis
port 389 nsew signal input
flabel metal2 s 440270 40710 440326 40910 0 FreeSans 320 90 0 0 gpio8_6_enable_inp_h
port 390 nsew signal input
flabel metal2 s 440856 40710 440908 40910 0 FreeSans 320 90 0 0 gpio8_6_enable_h
port 391 nsew signal input
flabel metal2 s 441585 40710 441637 40910 0 FreeSans 320 90 0 0 gpio8_6_hld_h_n
port 392 nsew signal input
flabel metal2 s 441899 40710 441951 40910 0 FreeSans 320 90 0 0 gpio8_6_analog_sel
port 393 nsew signal input
flabel metal2 s 442250 40710 442302 40910 0 FreeSans 320 90 0 0 gpio8_6_dm[2]
port 394 nsew signal input
flabel metal2 s 434581 40710 434633 40910 0 FreeSans 320 90 0 0 gpio8_6_dm[1]
port 395 nsew signal input
flabel metal2 s 437977 40710 438029 40910 0 FreeSans 320 90 0 0 gpio8_6_dm[0]
port 396 nsew signal input
flabel metal2 s 442628 40710 442680 40910 0 FreeSans 320 90 0 0 gpio8_6_hld_ovr
port 397 nsew signal input
flabel metal2 s 443477 40710 443529 40910 0 FreeSans 320 90 0 0 gpio8_6_out
port 398 nsew signal input
flabel metal2 s 444686 40710 444738 40910 0 FreeSans 320 90 0 0 gpio8_6_enable_vswitch_h
port 399 nsew signal input
flabel metal2 s 445397 40710 445449 40910 0 FreeSans 320 90 0 0 gpio8_6_enable_vdda_h
port 400 nsew signal input
flabel metal2 s 446645 40710 446697 40910 0 FreeSans 320 90 0 0 gpio8_6_vtrip_sel
port 401 nsew signal input
flabel metal2 s 446965 40710 447017 40910 0 FreeSans 320 90 0 0 gpio8_6_ib_mode_sel
port 402 nsew signal input
flabel metal2 s 447279 40710 447331 40910 0 FreeSans 320 90 0 0 gpio8_6_oe_n
port 403 nsew signal input
flabel metal2 s 447797 40710 447921 40910 0 FreeSans 320 90 0 0 gpio8_6_in_h
port 404 nsew signal input
flabel metal2 s 430493 40710 430545 40910 0 FreeSans 320 90 0 0 gpio8_6_zero
port 405 nsew signal output
flabel metal2 s 430131 40710 430183 40910 0 FreeSans 320 90 0 0 gpio8_6_one
port 406 nsew signal output
flabel metal2 s 454457 40710 454509 40910 0 FreeSans 320 90 0 0 gpio8_7_tie_lo_esd
port 407 nsew signal output
flabel metal2 s 454757 40710 454809 40910 0 FreeSans 320 90 0 0 gpio8_7_in
port 408 nsew signal output
flabel metal2 s 455059 40710 455111 40910 0 FreeSans 320 90 0 0 gpio8_7_tie_hi_esd
port 409 nsew signal output
flabel metal2 s 455357 40710 455409 40910 0 FreeSans 320 90 0 0 gpio8_7_enable_vddio
port 410 nsew signal input
flabel metal2 s 455657 40710 455709 40910 0 FreeSans 320 90 0 0 gpio8_7_slow
port 411 nsew signal input
flabel metal2 s 455957 40710 456085 40910 0 FreeSans 320 90 0 0 gpio8_7_pad_a_esd_0_h
port 412 nsew signal bidirectional
flabel metal2 s 457215 40710 457345 40910 0 FreeSans 320 90 0 0 gpio8_7_pad_a_esd_1_h
port 413 nsew signal bidirectional
flabel metal2 s 458223 40710 458437 40910 0 FreeSans 320 90 0 0 gpio8_7_pad_a_noesd_h
port 414 nsew signal bidirectional
flabel metal2 s 458689 40710 458741 40910 0 FreeSans 320 90 0 0 gpio8_7_analog_en
port 415 nsew signal input
flabel metal2 s 461603 40710 461655 40910 0 FreeSans 320 90 0 0 gpio8_7_analog_pol
port 416 nsew signal input
flabel metal2 s 461899 40710 461951 40910 0 FreeSans 320 90 0 0 gpio8_7_inp_dis
port 417 nsew signal input
flabel metal2 s 463270 40710 463326 40910 0 FreeSans 320 90 0 0 gpio8_7_enable_inp_h
port 418 nsew signal input
flabel metal2 s 463856 40710 463908 40910 0 FreeSans 320 90 0 0 gpio8_7_enable_h
port 419 nsew signal input
flabel metal2 s 464585 40710 464637 40910 0 FreeSans 320 90 0 0 gpio8_7_hld_h_n
port 420 nsew signal input
flabel metal2 s 464899 40710 464951 40910 0 FreeSans 320 90 0 0 gpio8_7_analog_sel
port 421 nsew signal input
flabel metal2 s 465250 40710 465302 40910 0 FreeSans 320 90 0 0 gpio8_7_dm[2]
port 422 nsew signal input
flabel metal2 s 457581 40710 457633 40910 0 FreeSans 320 90 0 0 gpio8_7_dm[1]
port 423 nsew signal input
flabel metal2 s 460977 40710 461029 40910 0 FreeSans 320 90 0 0 gpio8_7_dm[0]
port 424 nsew signal input
flabel metal2 s 465628 40710 465680 40910 0 FreeSans 320 90 0 0 gpio8_7_hld_ovr
port 425 nsew signal input
flabel metal2 s 466477 40710 466529 40910 0 FreeSans 320 90 0 0 gpio8_7_out
port 426 nsew signal input
flabel metal2 s 467686 40710 467738 40910 0 FreeSans 320 90 0 0 gpio8_7_enable_vswitch_h
port 427 nsew signal input
flabel metal2 s 468397 40710 468449 40910 0 FreeSans 320 90 0 0 gpio8_7_enable_vdda_h
port 428 nsew signal input
flabel metal2 s 469645 40710 469697 40910 0 FreeSans 320 90 0 0 gpio8_7_vtrip_sel
port 429 nsew signal input
flabel metal2 s 469965 40710 470017 40910 0 FreeSans 320 90 0 0 gpio8_7_ib_mode_sel
port 430 nsew signal input
flabel metal2 s 470279 40710 470331 40910 0 FreeSans 320 90 0 0 gpio8_7_oe_n
port 431 nsew signal input
flabel metal2 s 470797 40710 470921 40910 0 FreeSans 320 90 0 0 gpio8_7_in_h
port 432 nsew signal input
flabel metal2 s 453493 40710 453545 40910 0 FreeSans 320 90 0 0 gpio8_7_zero
port 433 nsew signal output
flabel metal2 s 453131 40710 453183 40910 0 FreeSans 320 90 0 0 gpio8_7_one
port 434 nsew signal output
flabel metal2 s 515865 40300 515917 40600 0 FreeSans 320 90 0 0 pwrdet_out2_vddio_hv
port 435 nsew signal output
flabel metal2 s 516097 40300 516149 40600 0 FreeSans 320 90 0 0 pwrdet_out1_vddd_hv
port 436 nsew signal output
flabel metal2 s 516344 40300 516396 40600 0 FreeSans 320 90 0 0 pwrdet_in1_vddio_hv
port 437 nsew signal input
flabel metal2 s 516556 40300 516608 40600 0 FreeSans 320 90 0 0 pwrdet_in2_vddd_hv
port 438 nsew signal input
flabel metal2 s 516896 40300 516948 40600 0 FreeSans 320 90 0 0 pwrdet_in1_vddd_hv
port 439 nsew signal input
flabel metal2 s 517210 40300 517262 40600 0 FreeSans 320 90 0 0 pwrdet_out1_vddio_hv
port 440 nsew signal output
flabel metal2 s 517427 40300 517479 40600 0 FreeSans 320 90 0 0 pwrdet_out2_vddd_hv
port 441 nsew signal output
flabel metal2 s 517659 40300 517711 40600 0 FreeSans 320 90 0 0 pwrdet_out3_vddd_hv
port 442 nsew signal output
flabel metal2 s 517952 40300 518004 40600 0 FreeSans 320 90 0 0 pwrdet_vddio_present_vddd_hv
port 443 nsew signal output
flabel metal2 s 519285 40300 519337 40600 0 FreeSans 320 90 0 0 pwrdet_out3_vddio_hv
port 444 nsew signal output
flabel metal2 s 523619 40300 523697 40600 0 FreeSans 320 90 0 0 pwrdet_tie_lo_esd
port 445 nsew signal output
flabel metal2 s 523965 40300 524017 40600 0 FreeSans 320 90 0 0 pwrdet_in3_vddd_hv
port 446 nsew signal input
flabel metal2 s 524219 40300 524271 40600 0 FreeSans 320 90 0 0 pwrdet_vddd_present_vddio_hv
port 447 nsew signal output
flabel metal2 s 524476 40300 524528 40600 0 FreeSans 320 90 0 0 pwrdet_in2_vddio_hv
port 448 nsew signal input
flabel metal2 s 524713 40300 524765 40600 0 FreeSans 320 90 0 0 pwrdet_in3_vddio_hv
port 449 nsew signal input
flabel metal2 s 525846 40300 525898 40600 0 FreeSans 320 90 0 0 pwrdet_rst_por_hv_n
port 450 nsew signal input
flabel metal2 s 576666 51043 576794 51343 0 FreeSans 320 90 0 0 sio_vinref_dft
port 451 nsew signal input
flabel metal2 s 576966 51043 577094 51343 0 FreeSans 320 90 0 0 sio_voutref_dft
port 452 nsew signal input
flabel metal2 s 579167 51043 579219 51343 0 FreeSans 320 90 0 0 sio_vref_sel[1]
port 453 nsew signal input
flabel metal2 s 579317 51043 579369 51343 0 FreeSans 320 90 0 0 sio_vref_sel[0]
port 454 nsew signal input
flabel metal2 s 579467 51043 579519 51343 0 FreeSans 320 90 0 0 sio_enable_vdda_h
port 455 nsew signal input
flabel metal2 s 579617 51043 579669 51343 0 FreeSans 320 90 0 0 sio_dft_refgen
port 456 nsew signal input
flabel metal2 s 579772 51043 579814 51343 0 FreeSans 320 90 0 0 sio_voh_sel[2]
port 457 nsew signal input
flabel metal2 s 579926 51043 579962 51343 0 FreeSans 320 90 0 0 sio_voh_sel[1]
port 458 nsew signal input
flabel metal2 s 580073 51043 580116 51343 0 FreeSans 320 90 0 0 sio_voh_sel[0]
port 459 nsew signal input
flabel metal2 s 368752 996600 368880 996900 0 FreeSans 320 90 0 0 amuxbus_a_n
port 460 nsew signal bidirectional
flabel metal2 s 368496 996600 368624 996900 0 FreeSans 320 90 0 0 amuxbus_b_n
port 461 nsew signal bidirectional
flabel metal2 s 580217 51043 580269 51343 0 FreeSans 320 90 0 0 sio_amuxbus_b
port 462 nsew analog bidirectional
flabel metal2 s 580367 51043 580419 51343 0 FreeSans 320 90 0 0 sio_amuxbus_a
port 463 nsew analog bidirectional
flabel metal2 s 580980 51043 581032 51343 0 FreeSans 320 90 0 0 sio_vreg_en_refgen
port 464 nsew signal input
flabel metal2 s 585410 51043 585462 51343 0 FreeSans 320 90 0 0 sio_ibuf_sel_refgen
port 465 nsew signal input
flabel metal2 s 586059 51043 586111 51343 0 FreeSans 320 90 0 0 sio_vohref
port 466 nsew signal input
flabel metal2 s 588949 51043 589001 51343 0 FreeSans 320 90 0 0 sio_hld_h_n_refgen
port 467 nsew signal input
flabel metal2 s 589380 51043 589432 51343 0 FreeSans 320 90 0 0 sio_vtrip_sel_refgen
port 468 nsew signal input
flabel metal2 s 609051 51043 609220 51343 0 FreeSans 320 90 0 0 sio_pad_a_esd_0_h[1]
port 469 nsew signal input
flabel metal2 s 609249 51043 609418 51343 0 FreeSans 320 90 0 0 sio_pad_a_noesd_h[1]
port 470 nsew signal input
flabel metal2 s 613341 51043 613393 51343 0 FreeSans 320 90 0 0 sio_inp_dis[1]
port 471 nsew signal input
flabel metal2 s 614017 51043 614069 51343 0 FreeSans 320 90 0 0 sio_tie_lo_esd[1]
port 472 nsew signal output
flabel metal2 s 616290 51043 616342 51343 0 FreeSans 320 90 0 0 sio_out[1]
port 473 nsew signal input
flabel metal2 s 617624 51043 617676 51343 0 FreeSans 320 90 0 0 sio_vtrip_sel[1]
port 474 nsew signal input
flabel metal2 s 619034 51043 619086 51343 0 FreeSans 320 90 0 0 sio_ibuf_sel[1]
port 475 nsew signal input
flabel metal2 s 619114 51043 619166 51343 0 FreeSans 320 90 0 0 sio_hld_h_n[1]
port 476 nsew signal input
flabel metal2 s 620239 51043 620308 51343 0 FreeSans 320 90 0 0 sio_hld_ovr[1]
port 477 nsew signal input
flabel metal2 s 620400 51043 620452 51343 0 FreeSans 320 90 0 0 sio_in[1]
port 478 nsew signal output
flabel metal2 s 620480 51043 620532 51343 0 FreeSans 320 90 0 0 sio_in_h[1]
port 479 nsew signal output
flabel metal2 s 621442 51043 621494 51343 0 FreeSans 320 90 0 0 sio_oe_n[1]
port 480 nsew signal input
flabel metal2 s 621522 51043 621574 51343 0 FreeSans 320 90 0 0 sio_slow[1]
port 481 nsew signal input
flabel metal2 s 621960 51043 622012 51343 0 FreeSans 320 90 0 0 sio_vreg_en[1]
port 482 nsew signal input
flabel metal2 s 622681 51043 622733 51343 0 FreeSans 320 90 0 0 sio_enable_h
port 483 nsew signal input
flabel metal2 s 622761 51043 622813 51343 0 FreeSans 320 90 0 0 sio_dm1[2]
port 484 nsew signal input
flabel metal2 s 623195 51043 623247 51343 0 FreeSans 320 90 0 0 sio_dm1[1]
port 485 nsew signal input
flabel metal2 s 623275 51043 623327 51343 0 FreeSans 320 90 0 0 sio_dm1[0]
port 486 nsew signal input
flabel metal2 s 627397 51043 627797 51343 0 FreeSans 320 90 0 0 sio_pad_a_esd_1_h[1]
port 487 nsew signal bidirectional
flabel metal2 s 634202 51043 634602 51343 0 FreeSans 320 90 0 0 sio_pad_a_esd_1_h[0]
port 488 nsew signal bidirectional
flabel metal2 s 638672 51043 638724 51343 0 FreeSans 320 90 0 0 sio_dm0[0]
port 489 nsew signal input
flabel metal2 s 638752 51043 638804 51343 0 FreeSans 320 90 0 0 sio_dm0[1]
port 490 nsew signal input
flabel metal2 s 639186 51043 639238 51343 0 FreeSans 320 90 0 0 sio_dm0[2]
port 491 nsew signal input
flabel metal2 s 639987 51043 640039 51343 0 FreeSans 320 90 0 0 sio_vreg_en[0]
port 492 nsew signal input
flabel metal2 s 640425 51043 640477 51343 0 FreeSans 320 90 0 0 sio_slow[0]
port 493 nsew signal input
flabel metal2 s 640505 51043 640557 51343 0 FreeSans 320 90 0 0 sio_oe_n[0]
port 494 nsew signal input
flabel metal2 s 641467 51043 641519 51343 0 FreeSans 320 90 0 0 sio_in_h[0]
port 495 nsew signal input
flabel metal2 s 641547 51043 641599 51343 0 FreeSans 320 90 0 0 sio_in[0]
port 496 nsew signal input
flabel metal2 s 641691 51043 641760 51343 0 FreeSans 320 90 0 0 sio_hld_ovr[0]
port 497 nsew signal input
flabel metal2 s 642833 51043 642885 51343 0 FreeSans 320 90 0 0 sio_hld_h_n[0]
port 498 nsew signal input
flabel metal2 s 642913 51043 642965 51343 0 FreeSans 320 90 0 0 sio_ibuf_sel[0]
port 499 nsew signal input
flabel metal2 s 644323 51043 644375 51343 0 FreeSans 320 90 0 0 sio_vtrip_sel[0]
port 500 nsew signal input
flabel metal2 s 645657 51043 645709 51343 0 FreeSans 320 90 0 0 sio_out[0]
port 501 nsew signal input
flabel metal2 s 647930 51043 647982 51343 0 FreeSans 320 90 0 0 sio_tie_lo_esd[0]
port 502 nsew signal output
flabel metal2 s 648606 51043 648658 51343 0 FreeSans 320 90 0 0 sio_inp_dis[0]
port 503 nsew signal input
flabel metal2 s 652581 51043 652751 51343 0 FreeSans 320 90 0 0 sio_pad_a_noesd_h[0]
port 504 nsew signal bidirectional
flabel metal2 s 652779 51043 652948 51343 0 FreeSans 320 90 0 0 sio_pad_a_esd_0_h[0]
port 505 nsew signal bidirectional
flabel metal3 s 676700 42386 677000 42446 0 FreeSans 320 0 0 0 muxsplit_se_hld_vdda_h_n
port 506 nsew signal input
flabel metal3 s 676700 43266 677000 43326 0 FreeSans 320 0 0 0 muxsplit_se_enable_vdda_h
port 507 nsew signal input
flabel metal3 s 676700 46888 677000 46948 0 FreeSans 320 0 0 0 muxsplit_se_switch_aa_sl
port 508 nsew signal input
flabel metal3 s 676700 47140 677000 47200 0 FreeSans 320 0 0 0 muxsplit_se_switch_aa_s0
port 509 nsew signal input
flabel metal3 s 676700 47392 677000 47452 0 FreeSans 320 0 0 0 muxsplit_se_switch_bb_s0
port 510 nsew signal input
flabel metal3 s 676700 47644 677000 47704 0 FreeSans 320 0 0 0 muxsplit_se_switch_bb_sl
port 511 nsew signal input
flabel metal3 s 676700 47896 677000 47956 0 FreeSans 320 0 0 0 muxsplit_se_switch_bb_sr
port 512 nsew signal input
flabel metal3 s 676700 48232 677000 48292 0 FreeSans 320 0 0 0 muxsplit_se_switch_aa_sr
port 513 nsew signal input
flabel metal3 s 676758 73928 677058 73998 0 FreeSans 320 0 0 0 gpio0_0_tie_lo_esd
port 514 nsew signal output
flabel metal3 s 676762 74506 677062 74576 0 FreeSans 320 0 0 0 gpio0_0_in
port 515 nsew signal output
flabel metal3 s 676758 74226 677058 74296 0 FreeSans 320 0 0 0 gpio0_0_tie_hi_esd
port 516 nsew signal output
flabel metal3 s 676758 74818 677058 74888 0 FreeSans 320 0 0 0 gpio0_0_enable_vddio
port 517 nsew signal input
flabel metal3 s 676758 75092 677058 75162 0 FreeSans 320 0 0 0 gpio0_0_slow
port 518 nsew signal input
flabel metal3 s 676758 75382 677058 75510 0 FreeSans 320 0 0 0 gpio0_0_pad_a_esd_0_h
port 519 nsew signal bidirectional
flabel metal3 s 676758 76812 677058 76942 0 FreeSans 320 0 0 0 gpio0_0_pad_a_esd_1_h
port 520 nsew signal bidirectional
flabel metal3 s 676758 77822 677058 78036 0 FreeSans 320 0 0 0 gpio0_0_pad_a_noesd_h
port 521 nsew signal bidirectional
flabel metal3 s 676758 78598 677058 78668 0 FreeSans 320 0 0 0 gpio0_0_analog_en
port 522 nsew signal input
flabel metal3 s 676758 81358 677058 81428 0 FreeSans 320 0 0 0 gpio0_0_analog_pol
port 523 nsew signal input
flabel metal3 s 676758 81938 677058 82008 0 FreeSans 320 0 0 0 gpio0_0_inp_dis
port 524 nsew signal input
flabel metal3 s 676758 83104 677058 83174 0 FreeSans 320 0 0 0 gpio0_0_enable_inp_h
port 525 nsew signal input
flabel metal3 s 676758 83560 677058 83630 0 FreeSans 320 0 0 0 gpio0_0_enable_h
port 526 nsew signal input
flabel metal3 s 676758 84014 677058 84084 0 FreeSans 320 0 0 0 gpio0_0_hld_h_n
port 527 nsew signal input
flabel metal3 s 676758 84632 677058 84702 0 FreeSans 320 0 0 0 gpio0_0_analog_sel
port 528 nsew signal input
flabel metal3 s 676758 85076 677058 85146 0 FreeSans 320 0 0 0 gpio0_0_dm[2]
port 529 nsew signal input
flabel metal3 s 676758 77402 677058 77472 0 FreeSans 320 0 0 0 gpio0_0_dm[1]
port 530 nsew signal input
flabel metal3 s 676758 80810 677058 80880 0 FreeSans 320 0 0 0 gpio0_0_dm[0]
port 531 nsew signal input
flabel metal3 s 676758 85560 677058 85630 0 FreeSans 320 0 0 0 gpio0_0_hld_ovr
port 532 nsew signal input
flabel metal3 s 676758 86332 677058 86402 0 FreeSans 320 0 0 0 gpio0_0_out
port 533 nsew signal input
flabel metal3 s 676758 87532 677058 87602 0 FreeSans 320 0 0 0 gpio0_0_enable_vswitch_h
port 534 nsew signal input
flabel metal3 s 676758 88252 677058 88322 0 FreeSans 320 0 0 0 gpio0_0_enable_vdda_h
port 535 nsew signal input
flabel metal3 s 676758 89114 677058 89184 0 FreeSans 320 0 0 0 gpio0_0_vtrip_sel
port 536 nsew signal input
flabel metal3 s 676758 89458 677058 89528 0 FreeSans 320 0 0 0 gpio0_0_ib_mode_sel
port 537 nsew signal input
flabel metal3 s 676758 89868 677058 89938 0 FreeSans 320 0 0 0 gpio0_0_oe_n
port 538 nsew signal input
flabel metal3 s 676758 90396 677058 90520 0 FreeSans 320 0 0 0 gpio0_0_in_h
port 539 nsew signal output
flabel metal3 s 676758 72728 677058 72798 0 FreeSans 320 0 0 0 gpio0_0_zero
port 540 nsew signal output
flabel metal3 s 676758 72278 677058 72348 0 FreeSans 320 0 0 0 gpio0_0_one
port 541 nsew signal output
flabel metal3 s 676758 94928 677058 94998 0 FreeSans 320 0 0 0 gpio0_1_tie_lo_esd
port 542 nsew signal output
flabel metal3 s 676762 95506 677062 95576 0 FreeSans 320 0 0 0 gpio0_1_in
port 543 nsew signal output
flabel metal3 s 676758 95226 677058 95296 0 FreeSans 320 0 0 0 gpio0_1_tie_hi_esd
port 544 nsew signal output
flabel metal3 s 676758 95818 677058 95888 0 FreeSans 320 0 0 0 gpio0_1_enable_vddio
port 545 nsew signal input
flabel metal3 s 676758 96092 677058 96162 0 FreeSans 320 0 0 0 gpio0_1_slow
port 546 nsew signal input
flabel metal3 s 676758 96382 677058 96510 0 FreeSans 320 0 0 0 gpio0_1_pad_a_esd_0_h
port 547 nsew signal bidirectional
flabel metal3 s 676758 97812 677058 97942 0 FreeSans 320 0 0 0 gpio0_1_pad_a_esd_1_h
port 548 nsew signal bidirectional
flabel metal3 s 676758 98822 677058 99036 0 FreeSans 320 0 0 0 gpio0_1_pad_a_noesd_h
port 549 nsew signal bidirectional
flabel metal3 s 676758 99598 677058 99668 0 FreeSans 320 0 0 0 gpio0_1_analog_en
port 550 nsew signal input
flabel metal3 s 676758 102358 677058 102428 0 FreeSans 320 0 0 0 gpio0_1_analog_pol
port 551 nsew signal input
flabel metal3 s 676758 102938 677058 103008 0 FreeSans 320 0 0 0 gpio0_1_inp_dis
port 552 nsew signal input
flabel metal3 s 676758 104104 677058 104174 0 FreeSans 320 0 0 0 gpio0_1_enable_inp_h
port 553 nsew signal input
flabel metal3 s 676758 104560 677058 104630 0 FreeSans 320 0 0 0 gpio0_1_enable_h
port 554 nsew signal input
flabel metal3 s 676758 105014 677058 105084 0 FreeSans 320 0 0 0 gpio0_1_hld_h_n
port 555 nsew signal input
flabel metal3 s 676758 105632 677058 105702 0 FreeSans 320 0 0 0 gpio0_1_analog_sel
port 556 nsew signal input
flabel metal3 s 676758 106076 677058 106146 0 FreeSans 320 0 0 0 gpio0_1_dm[2]
port 557 nsew signal input
flabel metal3 s 676758 98402 677058 98472 0 FreeSans 320 0 0 0 gpio0_1_dm[1]
port 558 nsew signal input
flabel metal3 s 676758 101810 677058 101880 0 FreeSans 320 0 0 0 gpio0_1_dm[0]
port 559 nsew signal input
flabel metal3 s 676758 106560 677058 106630 0 FreeSans 320 0 0 0 gpio0_1_hld_ovr
port 560 nsew signal input
flabel metal3 s 676758 107332 677058 107402 0 FreeSans 320 0 0 0 gpio0_1_out
port 561 nsew signal input
flabel metal3 s 676758 108532 677058 108602 0 FreeSans 320 0 0 0 gpio0_1_enable_vswitch_h
port 562 nsew signal input
flabel metal3 s 676758 109252 677058 109322 0 FreeSans 320 0 0 0 gpio0_1_enable_vdda_h
port 563 nsew signal input
flabel metal3 s 676758 110114 677058 110184 0 FreeSans 320 0 0 0 gpio0_1_vtrip_sel
port 564 nsew signal input
flabel metal3 s 676758 110458 677058 110528 0 FreeSans 320 0 0 0 gpio0_1_ib_mode_sel
port 565 nsew signal input
flabel metal3 s 676758 110868 677058 110938 0 FreeSans 320 0 0 0 gpio0_1_oe_n
port 566 nsew signal input
flabel metal3 s 676758 111396 677058 111520 0 FreeSans 320 0 0 0 gpio0_1_in_h
port 567 nsew signal output
flabel metal3 s 676758 93728 677058 93798 0 FreeSans 320 0 0 0 gpio0_1_zero
port 568 nsew signal output
flabel metal3 s 676758 93278 677058 93348 0 FreeSans 320 0 0 0 gpio0_1_one
port 569 nsew signal output
flabel metal3 s 676758 115928 677058 115998 0 FreeSans 320 0 0 0 gpio0_2_tie_lo_esd
port 570 nsew signal output
flabel metal3 s 676762 116506 677062 116576 0 FreeSans 320 0 0 0 gpio0_2_in
port 571 nsew signal output
flabel metal3 s 676758 116226 677058 116296 0 FreeSans 320 0 0 0 gpio0_2_tie_hi_esd
port 572 nsew signal output
flabel metal3 s 676758 116818 677058 116888 0 FreeSans 320 0 0 0 gpio0_2_enable_vddio
port 573 nsew signal input
flabel metal3 s 676758 117092 677058 117162 0 FreeSans 320 0 0 0 gpio0_2_slow
port 574 nsew signal input
flabel metal3 s 676758 117382 677058 117510 0 FreeSans 320 0 0 0 gpio0_2_pad_a_esd_0_h
port 575 nsew signal bidirectional
flabel metal3 s 676758 118812 677058 118942 0 FreeSans 320 0 0 0 gpio0_2_pad_a_esd_1_h
port 576 nsew signal bidirectional
flabel metal3 s 676758 119822 677058 120036 0 FreeSans 320 0 0 0 gpio0_2_pad_a_noesd_h
port 577 nsew signal bidirectional
flabel metal3 s 676758 120598 677058 120668 0 FreeSans 320 0 0 0 gpio0_2_analog_en
port 578 nsew signal input
flabel metal3 s 676758 123358 677058 123428 0 FreeSans 320 0 0 0 gpio0_2_analog_pol
port 579 nsew signal input
flabel metal3 s 676758 123938 677058 124008 0 FreeSans 320 0 0 0 gpio0_2_inp_dis
port 580 nsew signal input
flabel metal3 s 676758 125104 677058 125174 0 FreeSans 320 0 0 0 gpio0_2_enable_inp_h
port 581 nsew signal input
flabel metal3 s 676758 125560 677058 125630 0 FreeSans 320 0 0 0 gpio0_2_enable_h
port 582 nsew signal input
flabel metal3 s 676758 126014 677058 126084 0 FreeSans 320 0 0 0 gpio0_2_hld_h_n
port 583 nsew signal input
flabel metal3 s 676758 126632 677058 126702 0 FreeSans 320 0 0 0 gpio0_2_analog_sel
port 584 nsew signal input
flabel metal3 s 676758 127076 677058 127146 0 FreeSans 320 0 0 0 gpio0_2_dm[2]
port 585 nsew signal input
flabel metal3 s 676758 119402 677058 119472 0 FreeSans 320 0 0 0 gpio0_2_dm[1]
port 586 nsew signal input
flabel metal3 s 676758 122810 677058 122880 0 FreeSans 320 0 0 0 gpio0_2_dm[0]
port 587 nsew signal input
flabel metal3 s 676758 127560 677058 127630 0 FreeSans 320 0 0 0 gpio0_2_hld_ovr
port 588 nsew signal input
flabel metal3 s 676758 128332 677058 128402 0 FreeSans 320 0 0 0 gpio0_2_out
port 589 nsew signal input
flabel metal3 s 676758 129532 677058 129602 0 FreeSans 320 0 0 0 gpio0_2_enable_vswitch_h
port 590 nsew signal input
flabel metal3 s 676758 130252 677058 130322 0 FreeSans 320 0 0 0 gpio0_2_enable_vdda_h
port 591 nsew signal input
flabel metal3 s 676758 131114 677058 131184 0 FreeSans 320 0 0 0 gpio0_2_vtrip_sel
port 592 nsew signal input
flabel metal3 s 676758 131458 677058 131528 0 FreeSans 320 0 0 0 gpio0_2_ib_mode_sel
port 593 nsew signal input
flabel metal3 s 676758 131868 677058 131938 0 FreeSans 320 0 0 0 gpio0_2_oe_n
port 594 nsew signal input
flabel metal3 s 676758 132396 677058 132520 0 FreeSans 320 0 0 0 gpio0_2_in_h
port 595 nsew signal output
flabel metal3 s 676758 114728 677058 114798 0 FreeSans 320 0 0 0 gpio0_2_zero
port 596 nsew signal output
flabel metal3 s 676758 114278 677058 114348 0 FreeSans 320 0 0 0 gpio0_2_one
port 597 nsew signal output
flabel metal3 s 676758 136928 677058 136998 0 FreeSans 320 0 0 0 gpio0_3_tie_lo_esd
port 598 nsew signal output
flabel metal3 s 676762 137506 677062 137576 0 FreeSans 320 0 0 0 gpio0_3_in
port 599 nsew signal output
flabel metal3 s 676758 137226 677058 137296 0 FreeSans 320 0 0 0 gpio0_3_tie_hi_esd
port 600 nsew signal output
flabel metal3 s 676758 137818 677058 137888 0 FreeSans 320 0 0 0 gpio0_3_enable_vddio
port 601 nsew signal input
flabel metal3 s 676758 138092 677058 138162 0 FreeSans 320 0 0 0 gpio0_3_slow
port 602 nsew signal input
flabel metal3 s 676758 138382 677058 138510 0 FreeSans 320 0 0 0 gpio0_3_pad_a_esd_0_h
port 603 nsew signal bidirectional
flabel metal3 s 676758 139812 677058 139942 0 FreeSans 320 0 0 0 gpio0_3_pad_a_esd_1_h
port 604 nsew signal bidirectional
flabel metal3 s 676758 140822 677058 141036 0 FreeSans 320 0 0 0 gpio0_3_pad_a_noesd_h
port 605 nsew signal bidirectional
flabel metal3 s 676758 141598 677058 141668 0 FreeSans 320 0 0 0 gpio0_3_analog_en
port 606 nsew signal input
flabel metal3 s 676758 144358 677058 144428 0 FreeSans 320 0 0 0 gpio0_3_analog_pol
port 607 nsew signal input
flabel metal3 s 676758 144938 677058 145008 0 FreeSans 320 0 0 0 gpio0_3_inp_dis
port 608 nsew signal input
flabel metal3 s 676758 146104 677058 146174 0 FreeSans 320 0 0 0 gpio0_3_enable_inp_h
port 609 nsew signal input
flabel metal3 s 676758 146560 677058 146630 0 FreeSans 320 0 0 0 gpio0_3_enable_h
port 610 nsew signal input
flabel metal3 s 676758 147014 677058 147084 0 FreeSans 320 0 0 0 gpio0_3_hld_h_n
port 611 nsew signal input
flabel metal3 s 676758 147632 677058 147702 0 FreeSans 320 0 0 0 gpio0_3_analog_sel
port 612 nsew signal input
flabel metal3 s 676758 148076 677058 148146 0 FreeSans 320 0 0 0 gpio0_3_dm[2]
port 613 nsew signal input
flabel metal3 s 676758 140402 677058 140472 0 FreeSans 320 0 0 0 gpio0_3_dm[1]
port 614 nsew signal input
flabel metal3 s 676758 143810 677058 143880 0 FreeSans 320 0 0 0 gpio0_3_dm[0]
port 615 nsew signal input
flabel metal3 s 676758 148560 677058 148630 0 FreeSans 320 0 0 0 gpio0_3_hld_ovr
port 616 nsew signal input
flabel metal3 s 676758 149332 677058 149402 0 FreeSans 320 0 0 0 gpio0_3_out
port 617 nsew signal input
flabel metal3 s 676758 150532 677058 150602 0 FreeSans 320 0 0 0 gpio0_3_enable_vswitch_h
port 618 nsew signal input
flabel metal3 s 676758 151252 677058 151322 0 FreeSans 320 0 0 0 gpio0_3_enable_vdda_h
port 619 nsew signal input
flabel metal3 s 676758 152114 677058 152184 0 FreeSans 320 0 0 0 gpio0_3_vtrip_sel
port 620 nsew signal input
flabel metal3 s 676758 152458 677058 152528 0 FreeSans 320 0 0 0 gpio0_3_ib_mode_sel
port 621 nsew signal input
flabel metal3 s 676758 152868 677058 152938 0 FreeSans 320 0 0 0 gpio0_3_oe_n
port 622 nsew signal input
flabel metal3 s 676758 153396 677058 153520 0 FreeSans 320 0 0 0 gpio0_3_in_h
port 623 nsew signal output
flabel metal3 s 676758 135728 677058 135798 0 FreeSans 320 0 0 0 gpio0_3_zero
port 624 nsew signal output
flabel metal3 s 676758 135278 677058 135348 0 FreeSans 320 0 0 0 gpio0_3_one
port 625 nsew signal output
flabel metal3 s 676758 197928 677058 197998 0 FreeSans 320 0 0 0 gpio0_4_tie_lo_esd
port 626 nsew signal output
flabel metal3 s 676762 198506 677062 198576 0 FreeSans 320 0 0 0 gpio0_4_in
port 627 nsew signal output
flabel metal3 s 676758 198226 677058 198296 0 FreeSans 320 0 0 0 gpio0_4_tie_hi_esd
port 628 nsew signal output
flabel metal3 s 676758 198818 677058 198888 0 FreeSans 320 0 0 0 gpio0_4_enable_vddio
port 629 nsew signal input
flabel metal3 s 676758 199092 677058 199162 0 FreeSans 320 0 0 0 gpio0_4_slow
port 630 nsew signal input
flabel metal3 s 676758 199382 677058 199510 0 FreeSans 320 0 0 0 gpio0_4_pad_a_esd_0_h
port 631 nsew signal bidirectional
flabel metal3 s 676758 200812 677058 200942 0 FreeSans 320 0 0 0 gpio0_4_pad_a_esd_1_h
port 632 nsew signal bidirectional
flabel metal3 s 676758 201822 677058 202036 0 FreeSans 320 0 0 0 gpio0_4_pad_a_noesd_h
port 633 nsew signal bidirectional
flabel metal3 s 676758 202598 677058 202668 0 FreeSans 320 0 0 0 gpio0_4_analog_en
port 634 nsew signal input
flabel metal3 s 676758 205358 677058 205428 0 FreeSans 320 0 0 0 gpio0_4_analog_pol
port 635 nsew signal input
flabel metal3 s 676758 205938 677058 206008 0 FreeSans 320 0 0 0 gpio0_4_inp_dis
port 636 nsew signal input
flabel metal3 s 676758 207104 677058 207174 0 FreeSans 320 0 0 0 gpio0_4_enable_inp_h
port 637 nsew signal input
flabel metal3 s 676758 207560 677058 207630 0 FreeSans 320 0 0 0 gpio0_4_enable_h
port 638 nsew signal input
flabel metal3 s 676758 208014 677058 208084 0 FreeSans 320 0 0 0 gpio0_4_hld_h_n
port 639 nsew signal input
flabel metal3 s 676758 208632 677058 208702 0 FreeSans 320 0 0 0 gpio0_4_analog_sel
port 640 nsew signal input
flabel metal3 s 676758 209076 677058 209146 0 FreeSans 320 0 0 0 gpio0_4_dm[2]
port 641 nsew signal input
flabel metal3 s 676758 201402 677058 201472 0 FreeSans 320 0 0 0 gpio0_4_dm[1]
port 642 nsew signal input
flabel metal3 s 676758 204810 677058 204880 0 FreeSans 320 0 0 0 gpio0_4_dm[0]
port 643 nsew signal input
flabel metal3 s 676758 209560 677058 209630 0 FreeSans 320 0 0 0 gpio0_4_hld_ovr
port 644 nsew signal input
flabel metal3 s 676758 210332 677058 210402 0 FreeSans 320 0 0 0 gpio0_4_out
port 645 nsew signal input
flabel metal3 s 676758 211532 677058 211602 0 FreeSans 320 0 0 0 gpio0_4_enable_vswitch_h
port 646 nsew signal input
flabel metal3 s 676758 212252 677058 212322 0 FreeSans 320 0 0 0 gpio0_4_enable_vdda_h
port 647 nsew signal input
flabel metal3 s 676758 213114 677058 213184 0 FreeSans 320 0 0 0 gpio0_4_vtrip_sel
port 648 nsew signal input
flabel metal3 s 676758 213458 677058 213528 0 FreeSans 320 0 0 0 gpio0_4_ib_mode_sel
port 649 nsew signal input
flabel metal3 s 676758 213868 677058 213938 0 FreeSans 320 0 0 0 gpio0_4_oe_n
port 650 nsew signal input
flabel metal3 s 676758 214396 677058 214520 0 FreeSans 320 0 0 0 gpio0_4_in_h
port 651 nsew signal output
flabel metal3 s 676758 196728 677058 196798 0 FreeSans 320 0 0 0 gpio0_4_zero
port 652 nsew signal output
flabel metal3 s 676758 196278 677058 196348 0 FreeSans 320 0 0 0 gpio0_4_one
port 653 nsew signal output
flabel metal3 s 676758 218928 677058 218998 0 FreeSans 320 0 0 0 gpio0_5_tie_lo_esd
port 654 nsew signal output
flabel metal3 s 676762 219506 677062 219576 0 FreeSans 320 0 0 0 gpio0_5_in
port 655 nsew signal output
flabel metal3 s 676758 219226 677058 219296 0 FreeSans 320 0 0 0 gpio0_5_tie_hi_esd
port 656 nsew signal output
flabel metal3 s 676758 219818 677058 219888 0 FreeSans 320 0 0 0 gpio0_5_enable_vddio
port 657 nsew signal input
flabel metal3 s 676758 220092 677058 220162 0 FreeSans 320 0 0 0 gpio0_5_slow
port 658 nsew signal input
flabel metal3 s 676758 220382 677058 220510 0 FreeSans 320 0 0 0 gpio0_5_pad_a_esd_0_h
port 659 nsew signal bidirectional
flabel metal3 s 676758 221812 677058 221942 0 FreeSans 320 0 0 0 gpio0_5_pad_a_esd_1_h
port 660 nsew signal bidirectional
flabel metal3 s 676758 222822 677058 223036 0 FreeSans 320 0 0 0 gpio0_5_pad_a_noesd_h
port 661 nsew signal bidirectional
flabel metal3 s 676758 223598 677058 223668 0 FreeSans 320 0 0 0 gpio0_5_analog_en
port 662 nsew signal input
flabel metal3 s 676758 226358 677058 226428 0 FreeSans 320 0 0 0 gpio0_5_analog_pol
port 663 nsew signal input
flabel metal3 s 676758 226938 677058 227008 0 FreeSans 320 0 0 0 gpio0_5_inp_dis
port 664 nsew signal input
flabel metal3 s 676758 228104 677058 228174 0 FreeSans 320 0 0 0 gpio0_5_enable_inp_h
port 665 nsew signal input
flabel metal3 s 676758 228560 677058 228630 0 FreeSans 320 0 0 0 gpio0_5_enable_h
port 666 nsew signal input
flabel metal3 s 676758 229014 677058 229084 0 FreeSans 320 0 0 0 gpio0_5_hld_h_n
port 667 nsew signal input
flabel metal3 s 676758 229632 677058 229702 0 FreeSans 320 0 0 0 gpio0_5_analog_sel
port 668 nsew signal input
flabel metal3 s 676758 230076 677058 230146 0 FreeSans 320 0 0 0 gpio0_5_dm[2]
port 669 nsew signal input
flabel metal3 s 676758 222402 677058 222472 0 FreeSans 320 0 0 0 gpio0_5_dm[1]
port 670 nsew signal input
flabel metal3 s 676758 225810 677058 225880 0 FreeSans 320 0 0 0 gpio0_5_dm[0]
port 671 nsew signal input
flabel metal3 s 676758 230560 677058 230630 0 FreeSans 320 0 0 0 gpio0_5_hld_ovr
port 672 nsew signal input
flabel metal3 s 676758 231332 677058 231402 0 FreeSans 320 0 0 0 gpio0_5_out
port 673 nsew signal input
flabel metal3 s 676758 232532 677058 232602 0 FreeSans 320 0 0 0 gpio0_5_enable_vswitch_h
port 674 nsew signal input
flabel metal3 s 676758 233252 677058 233322 0 FreeSans 320 0 0 0 gpio0_5_enable_vdda_h
port 675 nsew signal input
flabel metal3 s 676758 234114 677058 234184 0 FreeSans 320 0 0 0 gpio0_5_vtrip_sel
port 676 nsew signal input
flabel metal3 s 676758 234458 677058 234528 0 FreeSans 320 0 0 0 gpio0_5_ib_mode_sel
port 677 nsew signal input
flabel metal3 s 676758 234868 677058 234938 0 FreeSans 320 0 0 0 gpio0_5_oe_n
port 678 nsew signal input
flabel metal3 s 676758 235396 677058 235520 0 FreeSans 320 0 0 0 gpio0_5_in_h
port 679 nsew signal output
flabel metal3 s 676758 217728 677058 217798 0 FreeSans 320 0 0 0 gpio0_5_zero
port 680 nsew signal output
flabel metal3 s 676758 217278 677058 217348 0 FreeSans 320 0 0 0 gpio0_5_one
port 681 nsew signal output
flabel metal3 s 676758 239928 677058 239998 0 FreeSans 320 0 0 0 gpio0_6_tie_lo_esd
port 682 nsew signal output
flabel metal3 s 676762 240506 677062 240576 0 FreeSans 320 0 0 0 gpio0_6_in
port 683 nsew signal output
flabel metal3 s 676758 240226 677058 240296 0 FreeSans 320 0 0 0 gpio0_6_tie_hi_esd
port 684 nsew signal output
flabel metal3 s 676758 240818 677058 240888 0 FreeSans 320 0 0 0 gpio0_6_enable_vddio
port 685 nsew signal input
flabel metal3 s 676758 241092 677058 241162 0 FreeSans 320 0 0 0 gpio0_6_slow
port 686 nsew signal input
flabel metal3 s 676758 241382 677058 241510 0 FreeSans 320 0 0 0 gpio0_6_pad_a_esd_0_h
port 687 nsew signal bidirectional
flabel metal3 s 676758 242812 677058 242942 0 FreeSans 320 0 0 0 gpio0_6_pad_a_esd_1_h
port 688 nsew signal bidirectional
flabel metal3 s 676758 243822 677058 244036 0 FreeSans 320 0 0 0 gpio0_6_pad_a_noesd_h
port 689 nsew signal bidirectional
flabel metal3 s 676758 244598 677058 244668 0 FreeSans 320 0 0 0 gpio0_6_analog_en
port 690 nsew signal input
flabel metal3 s 676758 247358 677058 247428 0 FreeSans 320 0 0 0 gpio0_6_analog_pol
port 691 nsew signal input
flabel metal3 s 676758 247938 677058 248008 0 FreeSans 320 0 0 0 gpio0_6_inp_dis
port 692 nsew signal input
flabel metal3 s 676758 249104 677058 249174 0 FreeSans 320 0 0 0 gpio0_6_enable_inp_h
port 693 nsew signal input
flabel metal3 s 676758 249560 677058 249630 0 FreeSans 320 0 0 0 gpio0_6_enable_h
port 694 nsew signal input
flabel metal3 s 676758 250014 677058 250084 0 FreeSans 320 0 0 0 gpio0_6_hld_h_n
port 695 nsew signal input
flabel metal3 s 676758 250632 677058 250702 0 FreeSans 320 0 0 0 gpio0_6_analog_sel
port 696 nsew signal input
flabel metal3 s 676758 251076 677058 251146 0 FreeSans 320 0 0 0 gpio0_6_dm[2]
port 697 nsew signal input
flabel metal3 s 676758 243402 677058 243472 0 FreeSans 320 0 0 0 gpio0_6_dm[1]
port 698 nsew signal input
flabel metal3 s 676758 246810 677058 246880 0 FreeSans 320 0 0 0 gpio0_6_dm[0]
port 699 nsew signal input
flabel metal3 s 676758 251560 677058 251630 0 FreeSans 320 0 0 0 gpio0_6_hld_ovr
port 700 nsew signal input
flabel metal3 s 676758 252332 677058 252402 0 FreeSans 320 0 0 0 gpio0_6_out
port 701 nsew signal input
flabel metal3 s 676758 253532 677058 253602 0 FreeSans 320 0 0 0 gpio0_6_enable_vswitch_h
port 702 nsew signal input
flabel metal3 s 676758 254252 677058 254322 0 FreeSans 320 0 0 0 gpio0_6_enable_vdda_h
port 703 nsew signal input
flabel metal3 s 676758 255114 677058 255184 0 FreeSans 320 0 0 0 gpio0_6_vtrip_sel
port 704 nsew signal input
flabel metal3 s 676758 255458 677058 255528 0 FreeSans 320 0 0 0 gpio0_6_ib_mode_sel
port 705 nsew signal input
flabel metal3 s 676758 255868 677058 255938 0 FreeSans 320 0 0 0 gpio0_6_oe_n
port 706 nsew signal input
flabel metal3 s 676758 256396 677058 256520 0 FreeSans 320 0 0 0 gpio0_6_in_h
port 707 nsew signal output
flabel metal3 s 676758 238728 677058 238798 0 FreeSans 320 0 0 0 gpio0_6_zero
port 708 nsew signal output
flabel metal3 s 676758 238278 677058 238348 0 FreeSans 320 0 0 0 gpio0_6_one
port 709 nsew signal output
flabel metal3 s 676758 260928 677058 260998 0 FreeSans 320 0 0 0 gpio0_7_tie_lo_esd
port 710 nsew signal output
flabel metal3 s 676762 261506 677062 261576 0 FreeSans 320 0 0 0 gpio0_7_in
port 711 nsew signal output
flabel metal3 s 676758 261226 677058 261296 0 FreeSans 320 0 0 0 gpio0_7_tie_hi_esd
port 712 nsew signal output
flabel metal3 s 676758 261818 677058 261888 0 FreeSans 320 0 0 0 gpio0_7_enable_vddio
port 713 nsew signal input
flabel metal3 s 676758 262092 677058 262162 0 FreeSans 320 0 0 0 gpio0_7_slow
port 714 nsew signal input
flabel metal3 s 676758 262382 677058 262510 0 FreeSans 320 0 0 0 gpio0_7_pad_a_esd_0_h
port 715 nsew signal bidirectional
flabel metal3 s 676758 263812 677058 263942 0 FreeSans 320 0 0 0 gpio0_7_pad_a_esd_1_h
port 716 nsew signal bidirectional
flabel metal3 s 676758 264822 677058 265036 0 FreeSans 320 0 0 0 gpio0_7_pad_a_noesd_h
port 717 nsew signal bidirectional
flabel metal3 s 676758 265598 677058 265668 0 FreeSans 320 0 0 0 gpio0_7_analog_en
port 718 nsew signal input
flabel metal3 s 676758 268358 677058 268428 0 FreeSans 320 0 0 0 gpio0_7_analog_pol
port 719 nsew signal input
flabel metal3 s 676758 268938 677058 269008 0 FreeSans 320 0 0 0 gpio0_7_inp_dis
port 720 nsew signal input
flabel metal3 s 676758 270104 677058 270174 0 FreeSans 320 0 0 0 gpio0_7_enable_inp_h
port 721 nsew signal input
flabel metal3 s 676758 270560 677058 270630 0 FreeSans 320 0 0 0 gpio0_7_enable_h
port 722 nsew signal input
flabel metal3 s 676758 271014 677058 271084 0 FreeSans 320 0 0 0 gpio0_7_hld_h_n
port 723 nsew signal input
flabel metal3 s 676758 271632 677058 271702 0 FreeSans 320 0 0 0 gpio0_7_analog_sel
port 724 nsew signal input
flabel metal3 s 676758 272076 677058 272146 0 FreeSans 320 0 0 0 gpio0_7_dm[2]
port 725 nsew signal input
flabel metal3 s 676758 264402 677058 264472 0 FreeSans 320 0 0 0 gpio0_7_dm[1]
port 726 nsew signal input
flabel metal3 s 676758 267810 677058 267880 0 FreeSans 320 0 0 0 gpio0_7_dm[0]
port 727 nsew signal input
flabel metal3 s 676758 272560 677058 272630 0 FreeSans 320 0 0 0 gpio0_7_hld_ovr
port 728 nsew signal input
flabel metal3 s 676758 273332 677058 273402 0 FreeSans 320 0 0 0 gpio0_7_out
port 729 nsew signal input
flabel metal3 s 676758 274532 677058 274602 0 FreeSans 320 0 0 0 gpio0_7_enable_vswitch_h
port 730 nsew signal input
flabel metal3 s 676758 275252 677058 275322 0 FreeSans 320 0 0 0 gpio0_7_enable_vdda_h
port 731 nsew signal input
flabel metal3 s 676758 276114 677058 276184 0 FreeSans 320 0 0 0 gpio0_7_vtrip_sel
port 732 nsew signal input
flabel metal3 s 676758 276458 677058 276528 0 FreeSans 320 0 0 0 gpio0_7_ib_mode_sel
port 733 nsew signal input
flabel metal3 s 676758 276868 677058 276938 0 FreeSans 320 0 0 0 gpio0_7_oe_n
port 734 nsew signal input
flabel metal3 s 676758 277396 677058 277520 0 FreeSans 320 0 0 0 gpio0_7_in_h
port 735 nsew signal output
flabel metal3 s 676758 259728 677058 259798 0 FreeSans 320 0 0 0 gpio0_7_zero
port 736 nsew signal output
flabel metal3 s 676758 259278 677058 259348 0 FreeSans 320 0 0 0 gpio0_7_one
port 737 nsew signal output
flabel metal3 s 677000 348539 677300 348605 0 FreeSans 320 0 0 0 gpio1_0_tie_hi_esd
port 738 nsew signal output
flabel metal3 s 677000 352855 677300 352921 0 FreeSans 320 0 0 0 gpio1_0_dm[2]
port 739 nsew signal input
flabel metal3 s 677000 348879 677300 348945 0 FreeSans 320 0 0 0 gpio1_0_dm[1]
port 740 nsew signal input
flabel metal3 s 677000 348709 677300 348775 0 FreeSans 320 0 0 0 gpio1_0_dm[0]
port 741 nsew signal input
flabel metal3 s 677000 349506 677300 349572 0 FreeSans 320 0 0 0 gpio1_0_slow
port 742 nsew signal input
flabel metal3 s 677000 349645 677300 349711 0 FreeSans 320 0 0 0 gpio1_0_oe_n
port 743 nsew signal input
flabel metal3 s 677000 351422 677300 351542 0 FreeSans 320 0 0 0 gpio1_0_tie_lo_esd
port 744 nsew signal output
flabel metal3 s 677000 353025 677300 353091 0 FreeSans 320 0 0 0 gpio1_0_inp_dis
port 745 nsew signal input
flabel metal3 s 677000 355357 677300 355431 0 FreeSans 320 0 0 0 gpio1_0_enable_vddio
port 746 nsew signal input
flabel metal3 s 677000 357001 677300 357067 0 FreeSans 320 0 0 0 gpio1_0_vtrip_sel
port 747 nsew signal input
flabel metal3 s 677000 361147 677300 361213 0 FreeSans 320 0 0 0 gpio1_0_ib_mode_sel[1]
port 748 nsew signal input
flabel metal3 s 677000 357171 677300 357237 0 FreeSans 320 0 0 0 gpio1_0_ib_mode_sel[0]
port 749 nsew signal input
flabel metal3 s 677000 359709 677300 359775 0 FreeSans 320 0 0 0 gpio1_0_out
port 750 nsew signal input
flabel metal3 s 677000 365293 677300 365359 0 FreeSans 320 0 0 0 gpio1_0_slew_ctl[1]
port 751 nsew signal input
flabel metal3 s 677000 361317 677300 361383 0 FreeSans 320 0 0 0 gpio1_0_slew_ctl[0]
port 752 nsew signal input
flabel metal3 s 677000 361487 677300 361553 0 FreeSans 320 0 0 0 gpio1_0_analog_pol
port 753 nsew signal input
flabel metal3 s 677000 364203 677300 364269 0 FreeSans 320 0 0 0 gpio1_0_analog_sel
port 754 nsew signal input
flabel metal3 s 677000 365463 677300 365529 0 FreeSans 320 0 0 0 gpio1_0_hys_trim
port 755 nsew signal input
flabel metal3 s 677000 365727 677300 365793 0 FreeSans 320 0 0 0 gpio1_0_vinref
port 756 nsew signal input
flabel metal3 s 677000 369063 677300 369129 0 FreeSans 320 0 0 0 gpio1_0_hld_ovr
port 757 nsew signal input
flabel metal3 s 677000 369658 677300 369724 0 FreeSans 320 0 0 0 gpio1_0_in_h
port 758 nsew signal output
flabel metal3 s 677000 370107 677300 370173 0 FreeSans 320 0 0 0 gpio1_0_enable_h
port 759 nsew signal input
flabel metal3 s 677000 370458 677300 370524 0 FreeSans 320 0 0 0 gpio1_0_in
port 760 nsew signal output
flabel metal3 s 677000 370607 677300 370673 0 FreeSans 320 0 0 0 gpio1_0_hld_h_n
port 761 nsew signal input
flabel metal3 s 677000 372780 677300 372846 0 FreeSans 320 0 0 0 gpio1_0_enable_vdda_h
port 762 nsew signal input
flabel metal3 s 677000 372911 677300 372977 0 FreeSans 320 0 0 0 gpio1_0_analog_en
port 763 nsew signal input
flabel metal3 s 677000 373112 677300 373178 0 FreeSans 320 0 0 0 gpio1_0_enable_inp_h
port 764 nsew signal input
flabel metal3 s 677000 373327 677300 373447 0 FreeSans 320 0 0 0 gpio1_0_enable_vswitch_h
port 765 nsew signal input
flabel metal3 s 677000 373903 677300 374023 0 FreeSans 320 0 0 0 gpio1_0_pad_a_noesd_h
port 766 nsew signal bidirectional
flabel metal3 s 677000 374160 677300 374279 0 FreeSans 320 0 0 0 gpio1_0_pad_a_esd_0_h
port 767 nsew signal bidirectional
flabel metal3 s 677000 374414 677300 374534 0 FreeSans 320 0 0 0 gpio1_0_pad_a_esd_1_h
port 768 nsew signal bidirectional
flabel metal3 s 677000 344728 677300 344798 0 FreeSans 320 0 0 0 gpio1_0_zero
port 769 nsew signal output
flabel metal3 s 677000 344278 677300 344348 0 FreeSans 320 0 0 0 gpio1_0_one
port 770 nsew signal output
flabel metal3 s 677000 381539 677300 381605 0 FreeSans 320 0 0 0 gpio1_1_tie_hi_esd
port 771 nsew signal output
flabel metal3 s 677000 385855 677300 385921 0 FreeSans 320 0 0 0 gpio1_1_dm[2]
port 772 nsew signal input
flabel metal3 s 677000 381879 677300 381945 0 FreeSans 320 0 0 0 gpio1_1_dm[1]
port 773 nsew signal input
flabel metal3 s 677000 381709 677300 381775 0 FreeSans 320 0 0 0 gpio1_1_dm[0]
port 774 nsew signal input
flabel metal3 s 677000 382506 677300 382572 0 FreeSans 320 0 0 0 gpio1_1_slow
port 775 nsew signal input
flabel metal3 s 677000 382645 677300 382711 0 FreeSans 320 0 0 0 gpio1_1_oe_n
port 776 nsew signal input
flabel metal3 s 677000 384422 677300 384542 0 FreeSans 320 0 0 0 gpio1_1_tie_lo_esd
port 777 nsew signal output
flabel metal3 s 677000 386025 677300 386091 0 FreeSans 320 0 0 0 gpio1_1_inp_dis
port 778 nsew signal input
flabel metal3 s 677000 388357 677300 388431 0 FreeSans 320 0 0 0 gpio1_1_enable_vddio
port 779 nsew signal input
flabel metal3 s 677000 390001 677300 390067 0 FreeSans 320 0 0 0 gpio1_1_vtrip_sel
port 780 nsew signal input
flabel metal3 s 677000 394147 677300 394213 0 FreeSans 320 0 0 0 gpio1_1_ib_mode_sel[1]
port 781 nsew signal input
flabel metal3 s 677000 390171 677300 390237 0 FreeSans 320 0 0 0 gpio1_1_ib_mode_sel[0]
port 782 nsew signal input
flabel metal3 s 677000 392709 677300 392775 0 FreeSans 320 0 0 0 gpio1_1_out
port 783 nsew signal input
flabel metal3 s 677000 398293 677300 398359 0 FreeSans 320 0 0 0 gpio1_1_slew_ctl[1]
port 784 nsew signal input
flabel metal3 s 677000 394317 677300 394383 0 FreeSans 320 0 0 0 gpio1_1_slew_ctl[0]
port 785 nsew signal input
flabel metal3 s 677000 394487 677300 394553 0 FreeSans 320 0 0 0 gpio1_1_analog_pol
port 786 nsew signal input
flabel metal3 s 677000 397203 677300 397269 0 FreeSans 320 0 0 0 gpio1_1_analog_sel
port 787 nsew signal input
flabel metal3 s 677000 398463 677300 398529 0 FreeSans 320 0 0 0 gpio1_1_hys_trim
port 788 nsew signal input
flabel metal3 s 677000 398727 677300 398793 0 FreeSans 320 0 0 0 gpio1_1_vinref
port 789 nsew signal input
flabel metal3 s 677000 402063 677300 402129 0 FreeSans 320 0 0 0 gpio1_1_hld_ovr
port 790 nsew signal input
flabel metal3 s 677000 402658 677300 402724 0 FreeSans 320 0 0 0 gpio1_1_in_h
port 791 nsew signal output
flabel metal3 s 677000 403107 677300 403173 0 FreeSans 320 0 0 0 gpio1_1_enable_h
port 792 nsew signal input
flabel metal3 s 677000 403458 677300 403524 0 FreeSans 320 0 0 0 gpio1_1_in
port 793 nsew signal output
flabel metal3 s 677000 403607 677300 403673 0 FreeSans 320 0 0 0 gpio1_1_hld_h_n
port 794 nsew signal input
flabel metal3 s 677000 405780 677300 405846 0 FreeSans 320 0 0 0 gpio1_1_enable_vdda_h
port 795 nsew signal input
flabel metal3 s 677000 405911 677300 405977 0 FreeSans 320 0 0 0 gpio1_1_analog_en
port 796 nsew signal input
flabel metal3 s 677000 406112 677300 406178 0 FreeSans 320 0 0 0 gpio1_1_enable_inp_h
port 797 nsew signal input
flabel metal3 s 677000 406327 677300 406447 0 FreeSans 320 0 0 0 gpio1_1_enable_vswitch_h
port 798 nsew signal input
flabel metal3 s 677000 406903 677300 407023 0 FreeSans 320 0 0 0 gpio1_1_pad_a_noesd_h
port 799 nsew signal bidirectional
flabel metal3 s 677000 407160 677300 407279 0 FreeSans 320 0 0 0 gpio1_1_pad_a_esd_0_h
port 800 nsew signal bidirectional
flabel metal3 s 677000 407414 677300 407534 0 FreeSans 320 0 0 0 gpio1_1_pad_a_esd_1_h
port 801 nsew signal bidirectional
flabel metal3 s 677000 377728 677300 377798 0 FreeSans 320 0 0 0 gpio1_1_zero
port 802 nsew signal output
flabel metal3 s 677000 377278 677300 377348 0 FreeSans 320 0 0 0 gpio1_1_one
port 803 nsew signal output
flabel metal3 s 677000 414539 677300 414605 0 FreeSans 320 0 0 0 gpio1_2_tie_hi_esd
port 804 nsew signal output
flabel metal3 s 677000 418855 677300 418921 0 FreeSans 320 0 0 0 gpio1_2_dm[2]
port 805 nsew signal input
flabel metal3 s 677000 414879 677300 414945 0 FreeSans 320 0 0 0 gpio1_2_dm[1]
port 806 nsew signal input
flabel metal3 s 677000 414709 677300 414775 0 FreeSans 320 0 0 0 gpio1_2_dm[0]
port 807 nsew signal input
flabel metal3 s 677000 415506 677300 415572 0 FreeSans 320 0 0 0 gpio1_2_slow
port 808 nsew signal input
flabel metal3 s 677000 415645 677300 415711 0 FreeSans 320 0 0 0 gpio1_2_oe_n
port 809 nsew signal input
flabel metal3 s 677000 417422 677300 417542 0 FreeSans 320 0 0 0 gpio1_2_tie_lo_esd
port 810 nsew signal output
flabel metal3 s 677000 419025 677300 419091 0 FreeSans 320 0 0 0 gpio1_2_inp_dis
port 811 nsew signal input
flabel metal3 s 677000 421357 677300 421431 0 FreeSans 320 0 0 0 gpio1_2_enable_vddio
port 812 nsew signal input
flabel metal3 s 677000 423001 677300 423067 0 FreeSans 320 0 0 0 gpio1_2_vtrip_sel
port 813 nsew signal input
flabel metal3 s 677000 427147 677300 427213 0 FreeSans 320 0 0 0 gpio1_2_ib_mode_sel[1]
port 814 nsew signal input
flabel metal3 s 677000 423171 677300 423237 0 FreeSans 320 0 0 0 gpio1_2_ib_mode_sel[0]
port 815 nsew signal input
flabel metal3 s 677000 425709 677300 425775 0 FreeSans 320 0 0 0 gpio1_2_out
port 816 nsew signal input
flabel metal3 s 677000 431293 677300 431359 0 FreeSans 320 0 0 0 gpio1_2_slew_ctl[1]
port 817 nsew signal input
flabel metal3 s 677000 427317 677300 427383 0 FreeSans 320 0 0 0 gpio1_2_slew_ctl[0]
port 818 nsew signal input
flabel metal3 s 677000 427487 677300 427553 0 FreeSans 320 0 0 0 gpio1_2_analog_pol
port 819 nsew signal input
flabel metal3 s 677000 430203 677300 430269 0 FreeSans 320 0 0 0 gpio1_2_analog_sel
port 820 nsew signal input
flabel metal3 s 677000 431463 677300 431529 0 FreeSans 320 0 0 0 gpio1_2_hys_trim
port 821 nsew signal input
flabel metal3 s 677000 431727 677300 431793 0 FreeSans 320 0 0 0 gpio1_2_vinref
port 822 nsew signal input
flabel metal3 s 677000 435063 677300 435129 0 FreeSans 320 0 0 0 gpio1_2_hld_ovr
port 823 nsew signal input
flabel metal3 s 677000 435658 677300 435724 0 FreeSans 320 0 0 0 gpio1_2_in_h
port 824 nsew signal output
flabel metal3 s 677000 436107 677300 436173 0 FreeSans 320 0 0 0 gpio1_2_enable_h
port 825 nsew signal input
flabel metal3 s 677000 436458 677300 436524 0 FreeSans 320 0 0 0 gpio1_2_in
port 826 nsew signal output
flabel metal3 s 677000 436607 677300 436673 0 FreeSans 320 0 0 0 gpio1_2_hld_h_n
port 827 nsew signal input
flabel metal3 s 677000 438780 677300 438846 0 FreeSans 320 0 0 0 gpio1_2_enable_vdda_h
port 828 nsew signal input
flabel metal3 s 677000 438911 677300 438977 0 FreeSans 320 0 0 0 gpio1_2_analog_en
port 829 nsew signal input
flabel metal3 s 677000 439112 677300 439178 0 FreeSans 320 0 0 0 gpio1_2_enable_inp_h
port 830 nsew signal input
flabel metal3 s 677000 439327 677300 439447 0 FreeSans 320 0 0 0 gpio1_2_enable_vswitch_h
port 831 nsew signal input
flabel metal3 s 677000 439903 677300 440023 0 FreeSans 320 0 0 0 gpio1_2_pad_a_noesd_h
port 832 nsew signal bidirectional
flabel metal3 s 677000 440160 677300 440279 0 FreeSans 320 0 0 0 gpio1_2_pad_a_esd_0_h
port 833 nsew signal bidirectional
flabel metal3 s 677000 440414 677300 440534 0 FreeSans 320 0 0 0 gpio1_2_pad_a_esd_1_h
port 834 nsew signal bidirectional
flabel metal3 s 677000 410728 677300 410798 0 FreeSans 320 0 0 0 gpio1_2_zero
port 835 nsew signal output
flabel metal3 s 677000 410278 677300 410348 0 FreeSans 320 0 0 0 gpio1_2_one
port 836 nsew signal output
flabel metal3 s 677000 447539 677300 447605 0 FreeSans 320 0 0 0 gpio1_3_tie_hi_esd
port 837 nsew signal output
flabel metal3 s 677000 451855 677300 451921 0 FreeSans 320 0 0 0 gpio1_3_dm[2]
port 838 nsew signal input
flabel metal3 s 677000 447879 677300 447945 0 FreeSans 320 0 0 0 gpio1_3_dm[1]
port 839 nsew signal input
flabel metal3 s 677000 447709 677300 447775 0 FreeSans 320 0 0 0 gpio1_3_dm[0]
port 840 nsew signal input
flabel metal3 s 677000 448506 677300 448572 0 FreeSans 320 0 0 0 gpio1_3_slow
port 841 nsew signal input
flabel metal3 s 677000 448645 677300 448711 0 FreeSans 320 0 0 0 gpio1_3_oe_n
port 842 nsew signal input
flabel metal3 s 677000 450422 677300 450542 0 FreeSans 320 0 0 0 gpio1_3_tie_lo_esd
port 843 nsew signal output
flabel metal3 s 677000 452025 677300 452091 0 FreeSans 320 0 0 0 gpio1_3_inp_dis
port 844 nsew signal input
flabel metal3 s 677000 454357 677300 454431 0 FreeSans 320 0 0 0 gpio1_3_enable_vddio
port 845 nsew signal input
flabel metal3 s 677000 456001 677300 456067 0 FreeSans 320 0 0 0 gpio1_3_vtrip_sel
port 846 nsew signal input
flabel metal3 s 677000 460147 677300 460213 0 FreeSans 320 0 0 0 gpio1_3_ib_mode_sel[1]
port 847 nsew signal input
flabel metal3 s 677000 456171 677300 456237 0 FreeSans 320 0 0 0 gpio1_3_ib_mode_sel[0]
port 848 nsew signal input
flabel metal3 s 677000 458709 677300 458775 0 FreeSans 320 0 0 0 gpio1_3_out
port 849 nsew signal input
flabel metal3 s 677000 464293 677300 464359 0 FreeSans 320 0 0 0 gpio1_3_slew_ctl[1]
port 850 nsew signal input
flabel metal3 s 677000 460317 677300 460383 0 FreeSans 320 0 0 0 gpio1_3_slew_ctl[0]
port 851 nsew signal input
flabel metal3 s 677000 460487 677300 460553 0 FreeSans 320 0 0 0 gpio1_3_analog_pol
port 852 nsew signal input
flabel metal3 s 677000 463203 677300 463269 0 FreeSans 320 0 0 0 gpio1_3_analog_sel
port 853 nsew signal input
flabel metal3 s 677000 464463 677300 464529 0 FreeSans 320 0 0 0 gpio1_3_hys_trim
port 854 nsew signal input
flabel metal3 s 677000 464727 677300 464793 0 FreeSans 320 0 0 0 gpio1_3_vinref
port 855 nsew signal input
flabel metal3 s 677000 468063 677300 468129 0 FreeSans 320 0 0 0 gpio1_3_hld_ovr
port 856 nsew signal input
flabel metal3 s 677000 468658 677300 468724 0 FreeSans 320 0 0 0 gpio1_3_in_h
port 857 nsew signal output
flabel metal3 s 677000 469107 677300 469173 0 FreeSans 320 0 0 0 gpio1_3_enable_h
port 858 nsew signal input
flabel metal3 s 677000 469458 677300 469524 0 FreeSans 320 0 0 0 gpio1_3_in
port 859 nsew signal output
flabel metal3 s 677000 469607 677300 469673 0 FreeSans 320 0 0 0 gpio1_3_hld_h_n
port 860 nsew signal input
flabel metal3 s 677000 471780 677300 471846 0 FreeSans 320 0 0 0 gpio1_3_enable_vdda_h
port 861 nsew signal input
flabel metal3 s 677000 471911 677300 471977 0 FreeSans 320 0 0 0 gpio1_3_analog_en
port 862 nsew signal input
flabel metal3 s 677000 472112 677300 472178 0 FreeSans 320 0 0 0 gpio1_3_enable_inp_h
port 863 nsew signal input
flabel metal3 s 677000 472327 677300 472447 0 FreeSans 320 0 0 0 gpio1_3_enable_vswitch_h
port 864 nsew signal input
flabel metal3 s 677000 472903 677300 473023 0 FreeSans 320 0 0 0 gpio1_3_pad_a_noesd_h
port 865 nsew signal bidirectional
flabel metal3 s 677000 473160 677300 473279 0 FreeSans 320 0 0 0 gpio1_3_pad_a_esd_0_h
port 866 nsew signal bidirectional
flabel metal3 s 677000 473414 677300 473534 0 FreeSans 320 0 0 0 gpio1_3_pad_a_esd_1_h
port 867 nsew signal bidirectional
flabel metal3 s 677000 443728 677300 443798 0 FreeSans 320 0 0 0 gpio1_3_zero
port 868 nsew signal output
flabel metal3 s 677000 443278 677300 443348 0 FreeSans 320 0 0 0 gpio1_3_one
port 869 nsew signal output
flabel metal3 s 676700 501464 677000 501524 0 FreeSans 320 0 0 0 vref_e_ref_sel[1]
port 870 nsew signal input
flabel metal3 s 676700 502445 677000 502505 0 FreeSans 320 0 0 0 vref_e_ref_sel[0]
port 871 nsew signal input
flabel metal3 s 676700 506975 677000 507103 0 FreeSans 320 0 0 0 vref_e_vinref
port 872 nsew signal output
flabel metal3 s 676700 507799 677000 507859 0 FreeSans 320 0 0 0 vref_e_ref_sel[2]
port 873 nsew signal input
flabel metal3 s 676700 507997 677000 508057 0 FreeSans 320 0 0 0 vref_e_enable_h
port 874 nsew signal input
flabel metal3 s 676700 508197 677000 508257 0 FreeSans 320 0 0 0 vref_e_hld_h_n
port 875 nsew signal input
flabel metal3 s 676700 508485 677000 508545 0 FreeSans 320 0 0 0 vref_e_vrefgen_en
port 876 nsew signal input
flabel metal3 s 676700 513313 677000 513373 0 FreeSans 320 0 0 0 vref_e_ref_sel[4]
port 877 nsew signal input
flabel metal3 s 676700 513565 677000 513625 0 FreeSans 320 0 0 0 vref_e_ref_sel[3]
port 878 nsew signal input
flabel metal3 s 677000 516161 677300 516561 0 FreeSans 320 0 0 0 vcap_e_cpos
port 879 nsew signal input
flabel metal3 s 677000 545139 677300 545205 0 FreeSans 320 0 0 0 gpio1_4_tie_hi_esd
port 880 nsew signal output
flabel metal3 s 677000 549455 677300 549521 0 FreeSans 320 0 0 0 gpio1_4_dm[2]
port 881 nsew signal input
flabel metal3 s 677000 545479 677300 545545 0 FreeSans 320 0 0 0 gpio1_4_dm[1]
port 882 nsew signal input
flabel metal3 s 677000 545309 677300 545375 0 FreeSans 320 0 0 0 gpio1_4_dm[0]
port 883 nsew signal input
flabel metal3 s 677000 546106 677300 546172 0 FreeSans 320 0 0 0 gpio1_4_slow
port 884 nsew signal input
flabel metal3 s 677000 546245 677300 546311 0 FreeSans 320 0 0 0 gpio1_4_oe_n
port 885 nsew signal input
flabel metal3 s 677000 548022 677300 548142 0 FreeSans 320 0 0 0 gpio1_4_tie_lo_esd
port 886 nsew signal output
flabel metal3 s 677000 549625 677300 549691 0 FreeSans 320 0 0 0 gpio1_4_inp_dis
port 887 nsew signal input
flabel metal3 s 677000 551957 677300 552031 0 FreeSans 320 0 0 0 gpio1_4_enable_vddio
port 888 nsew signal input
flabel metal3 s 677000 553601 677300 553667 0 FreeSans 320 0 0 0 gpio1_4_vtrip_sel
port 889 nsew signal input
flabel metal3 s 677000 557747 677300 557813 0 FreeSans 320 0 0 0 gpio1_4_ib_mode_sel[1]
port 890 nsew signal input
flabel metal3 s 677000 553771 677300 553837 0 FreeSans 320 0 0 0 gpio1_4_ib_mode_sel[0]
port 891 nsew signal input
flabel metal3 s 677000 556309 677300 556375 0 FreeSans 320 0 0 0 gpio1_4_out
port 892 nsew signal input
flabel metal3 s 677000 561893 677300 561959 0 FreeSans 320 0 0 0 gpio1_4_slew_ctl[1]
port 893 nsew signal input
flabel metal3 s 677000 557917 677300 557983 0 FreeSans 320 0 0 0 gpio1_4_slew_ctl[0]
port 894 nsew signal input
flabel metal3 s 677000 558087 677300 558153 0 FreeSans 320 0 0 0 gpio1_4_analog_pol
port 895 nsew signal input
flabel metal3 s 677000 560803 677300 560869 0 FreeSans 320 0 0 0 gpio1_4_analog_sel
port 896 nsew signal input
flabel metal3 s 677000 562063 677300 562129 0 FreeSans 320 0 0 0 gpio1_4_hys_trim
port 897 nsew signal input
flabel metal3 s 677000 562327 677300 562393 0 FreeSans 320 0 0 0 gpio1_4_vinref
port 898 nsew signal input
flabel metal3 s 677000 565663 677300 565729 0 FreeSans 320 0 0 0 gpio1_4_hld_ovr
port 899 nsew signal input
flabel metal3 s 677000 566258 677300 566324 0 FreeSans 320 0 0 0 gpio1_4_in_h
port 900 nsew signal output
flabel metal3 s 677000 566707 677300 566773 0 FreeSans 320 0 0 0 gpio1_4_enable_h
port 901 nsew signal input
flabel metal3 s 677000 567058 677300 567124 0 FreeSans 320 0 0 0 gpio1_4_in
port 902 nsew signal output
flabel metal3 s 677000 567207 677300 567273 0 FreeSans 320 0 0 0 gpio1_4_hld_h_n
port 903 nsew signal input
flabel metal3 s 677000 569380 677300 569446 0 FreeSans 320 0 0 0 gpio1_4_enable_vdda_h
port 904 nsew signal input
flabel metal3 s 677000 569511 677300 569577 0 FreeSans 320 0 0 0 gpio1_4_analog_en
port 905 nsew signal input
flabel metal3 s 677000 569712 677300 569778 0 FreeSans 320 0 0 0 gpio1_4_enable_inp_h
port 906 nsew signal input
flabel metal3 s 677000 569927 677300 570047 0 FreeSans 320 0 0 0 gpio1_4_enable_vswitch_h
port 907 nsew signal input
flabel metal3 s 677000 570503 677300 570623 0 FreeSans 320 0 0 0 gpio1_4_pad_a_noesd_h
port 908 nsew signal bidirectional
flabel metal3 s 677000 570760 677300 570879 0 FreeSans 320 0 0 0 gpio1_4_pad_a_esd_0_h
port 909 nsew signal bidirectional
flabel metal3 s 677000 571014 677300 571134 0 FreeSans 320 0 0 0 gpio1_4_pad_a_esd_1_h
port 910 nsew signal bidirectional
flabel metal3 s 677000 541328 677300 541398 0 FreeSans 320 0 0 0 gpio1_4_zero
port 911 nsew signal output
flabel metal3 s 677000 540878 677300 540948 0 FreeSans 320 0 0 0 gpio1_4_one
port 912 nsew signal output
flabel metal3 s 677000 578139 677300 578205 0 FreeSans 320 0 0 0 gpio1_5_tie_hi_esd
port 913 nsew signal output
flabel metal3 s 677000 582455 677300 582521 0 FreeSans 320 0 0 0 gpio1_5_dm[2]
port 914 nsew signal input
flabel metal3 s 677000 578479 677300 578545 0 FreeSans 320 0 0 0 gpio1_5_dm[1]
port 915 nsew signal input
flabel metal3 s 677000 578309 677300 578375 0 FreeSans 320 0 0 0 gpio1_5_dm[0]
port 916 nsew signal input
flabel metal3 s 677000 579106 677300 579172 0 FreeSans 320 0 0 0 gpio1_5_slow
port 917 nsew signal input
flabel metal3 s 677000 579245 677300 579311 0 FreeSans 320 0 0 0 gpio1_5_oe_n
port 918 nsew signal input
flabel metal3 s 677000 581022 677300 581142 0 FreeSans 320 0 0 0 gpio1_5_tie_lo_esd
port 919 nsew signal output
flabel metal3 s 677000 582625 677300 582691 0 FreeSans 320 0 0 0 gpio1_5_inp_dis
port 920 nsew signal input
flabel metal3 s 677000 584957 677300 585031 0 FreeSans 320 0 0 0 gpio1_5_enable_vddio
port 921 nsew signal input
flabel metal3 s 677000 586601 677300 586667 0 FreeSans 320 0 0 0 gpio1_5_vtrip_sel
port 922 nsew signal input
flabel metal3 s 677000 590747 677300 590813 0 FreeSans 320 0 0 0 gpio1_5_ib_mode_sel[1]
port 923 nsew signal input
flabel metal3 s 677000 586771 677300 586837 0 FreeSans 320 0 0 0 gpio1_5_ib_mode_sel[0]
port 924 nsew signal input
flabel metal3 s 677000 589309 677300 589375 0 FreeSans 320 0 0 0 gpio1_5_out
port 925 nsew signal input
flabel metal3 s 677000 594893 677300 594959 0 FreeSans 320 0 0 0 gpio1_5_slew_ctl[1]
port 926 nsew signal input
flabel metal3 s 677000 590917 677300 590983 0 FreeSans 320 0 0 0 gpio1_5_slew_ctl[0]
port 927 nsew signal input
flabel metal3 s 677000 591087 677300 591153 0 FreeSans 320 0 0 0 gpio1_5_analog_pol
port 928 nsew signal input
flabel metal3 s 677000 593803 677300 593869 0 FreeSans 320 0 0 0 gpio1_5_analog_sel
port 929 nsew signal input
flabel metal3 s 677000 595063 677300 595129 0 FreeSans 320 0 0 0 gpio1_5_hys_trim
port 930 nsew signal input
flabel metal3 s 677000 595327 677300 595393 0 FreeSans 320 0 0 0 gpio1_5_vinref
port 931 nsew signal input
flabel metal3 s 677000 598663 677300 598729 0 FreeSans 320 0 0 0 gpio1_5_hld_ovr
port 932 nsew signal input
flabel metal3 s 677000 599258 677300 599324 0 FreeSans 320 0 0 0 gpio1_5_in_h
port 933 nsew signal output
flabel metal3 s 677000 599707 677300 599773 0 FreeSans 320 0 0 0 gpio1_5_enable_h
port 934 nsew signal input
flabel metal3 s 677000 600058 677300 600124 0 FreeSans 320 0 0 0 gpio1_5_in
port 935 nsew signal output
flabel metal3 s 677000 600207 677300 600273 0 FreeSans 320 0 0 0 gpio1_5_hld_h_n
port 936 nsew signal input
flabel metal3 s 677000 602380 677300 602446 0 FreeSans 320 0 0 0 gpio1_5_enable_vdda_h
port 937 nsew signal input
flabel metal3 s 677000 602511 677300 602577 0 FreeSans 320 0 0 0 gpio1_5_analog_en
port 938 nsew signal input
flabel metal3 s 677000 602712 677300 602778 0 FreeSans 320 0 0 0 gpio1_5_enable_inp_h
port 939 nsew signal input
flabel metal3 s 677000 602927 677300 603047 0 FreeSans 320 0 0 0 gpio1_5_enable_vswitch_h
port 940 nsew signal input
flabel metal3 s 677000 603503 677300 603623 0 FreeSans 320 0 0 0 gpio1_5_pad_a_noesd_h
port 941 nsew signal bidirectional
flabel metal3 s 677000 603760 677300 603879 0 FreeSans 320 0 0 0 gpio1_5_pad_a_esd_0_h
port 942 nsew signal bidirectional
flabel metal3 s 677000 604014 677300 604134 0 FreeSans 320 0 0 0 gpio1_5_pad_a_esd_1_h
port 943 nsew signal bidirectional
flabel metal3 s 677000 574328 677300 574398 0 FreeSans 320 0 0 0 gpio1_5_zero
port 944 nsew signal output
flabel metal3 s 677000 573878 677300 573948 0 FreeSans 320 0 0 0 gpio1_5_one
port 945 nsew signal output
flabel metal3 s 677000 611139 677300 611205 0 FreeSans 320 0 0 0 gpio1_6_tie_hi_esd
port 946 nsew signal output
flabel metal3 s 677000 615455 677300 615521 0 FreeSans 320 0 0 0 gpio1_6_dm[2]
port 947 nsew signal input
flabel metal3 s 677000 611479 677300 611545 0 FreeSans 320 0 0 0 gpio1_6_dm[1]
port 948 nsew signal input
flabel metal3 s 677000 611309 677300 611375 0 FreeSans 320 0 0 0 gpio1_6_dm[0]
port 949 nsew signal input
flabel metal3 s 677000 612106 677300 612172 0 FreeSans 320 0 0 0 gpio1_6_slow
port 950 nsew signal input
flabel metal3 s 677000 612245 677300 612311 0 FreeSans 320 0 0 0 gpio1_6_oe_n
port 951 nsew signal input
flabel metal3 s 677000 614022 677300 614142 0 FreeSans 320 0 0 0 gpio1_6_tie_lo_esd
port 952 nsew signal output
flabel metal3 s 677000 615625 677300 615691 0 FreeSans 320 0 0 0 gpio1_6_inp_dis
port 953 nsew signal input
flabel metal3 s 677000 617957 677300 618031 0 FreeSans 320 0 0 0 gpio1_6_enable_vddio
port 954 nsew signal input
flabel metal3 s 677000 619601 677300 619667 0 FreeSans 320 0 0 0 gpio1_6_vtrip_sel
port 955 nsew signal input
flabel metal3 s 677000 623747 677300 623813 0 FreeSans 320 0 0 0 gpio1_6_ib_mode_sel[1]
port 956 nsew signal input
flabel metal3 s 677000 619771 677300 619837 0 FreeSans 320 0 0 0 gpio1_6_ib_mode_sel[0]
port 957 nsew signal input
flabel metal3 s 677000 622309 677300 622375 0 FreeSans 320 0 0 0 gpio1_6_out
port 958 nsew signal input
flabel metal3 s 677000 627893 677300 627959 0 FreeSans 320 0 0 0 gpio1_6_slew_ctl[1]
port 959 nsew signal input
flabel metal3 s 677000 623917 677300 623983 0 FreeSans 320 0 0 0 gpio1_6_slew_ctl[0]
port 960 nsew signal input
flabel metal3 s 677000 624087 677300 624153 0 FreeSans 320 0 0 0 gpio1_6_analog_pol
port 961 nsew signal input
flabel metal3 s 677000 626803 677300 626869 0 FreeSans 320 0 0 0 gpio1_6_analog_sel
port 962 nsew signal input
flabel metal3 s 677000 628063 677300 628129 0 FreeSans 320 0 0 0 gpio1_6_hys_trim
port 963 nsew signal input
flabel metal3 s 677000 628327 677300 628393 0 FreeSans 320 0 0 0 gpio1_6_vinref
port 964 nsew signal input
flabel metal3 s 677000 631663 677300 631729 0 FreeSans 320 0 0 0 gpio1_6_hld_ovr
port 965 nsew signal input
flabel metal3 s 677000 632258 677300 632324 0 FreeSans 320 0 0 0 gpio1_6_in_h
port 966 nsew signal output
flabel metal3 s 677000 632707 677300 632773 0 FreeSans 320 0 0 0 gpio1_6_enable_h
port 967 nsew signal input
flabel metal3 s 677000 633058 677300 633124 0 FreeSans 320 0 0 0 gpio1_6_in
port 968 nsew signal output
flabel metal3 s 677000 633207 677300 633273 0 FreeSans 320 0 0 0 gpio1_6_hld_h_n
port 969 nsew signal input
flabel metal3 s 677000 635380 677300 635446 0 FreeSans 320 0 0 0 gpio1_6_enable_vdda_h
port 970 nsew signal input
flabel metal3 s 677000 635511 677300 635577 0 FreeSans 320 0 0 0 gpio1_6_analog_en
port 971 nsew signal input
flabel metal3 s 677000 635712 677300 635778 0 FreeSans 320 0 0 0 gpio1_6_enable_inp_h
port 972 nsew signal input
flabel metal3 s 677000 635927 677300 636047 0 FreeSans 320 0 0 0 gpio1_6_enable_vswitch_h
port 973 nsew signal input
flabel metal3 s 677000 636503 677300 636623 0 FreeSans 320 0 0 0 gpio1_6_pad_a_noesd_h
port 974 nsew signal bidirectional
flabel metal3 s 677000 636760 677300 636879 0 FreeSans 320 0 0 0 gpio1_6_pad_a_esd_0_h
port 975 nsew signal bidirectional
flabel metal3 s 677000 637014 677300 637134 0 FreeSans 320 0 0 0 gpio1_6_pad_a_esd_1_h
port 976 nsew signal bidirectional
flabel metal3 s 677000 607328 677300 607398 0 FreeSans 320 0 0 0 gpio1_6_zero
port 977 nsew signal output
flabel metal3 s 677000 606878 677300 606948 0 FreeSans 320 0 0 0 gpio1_6_one
port 978 nsew signal output
flabel metal3 s 677000 644139 677300 644205 0 FreeSans 320 0 0 0 gpio1_7_tie_hi_esd
port 979 nsew signal output
flabel metal3 s 677000 648455 677300 648521 0 FreeSans 320 0 0 0 gpio1_7_dm[2]
port 980 nsew signal input
flabel metal3 s 677000 644479 677300 644545 0 FreeSans 320 0 0 0 gpio1_7_dm[1]
port 981 nsew signal input
flabel metal3 s 677000 644309 677300 644375 0 FreeSans 320 0 0 0 gpio1_7_dm[0]
port 982 nsew signal input
flabel metal3 s 677000 645106 677300 645172 0 FreeSans 320 0 0 0 gpio1_7_slow
port 983 nsew signal input
flabel metal3 s 677000 645245 677300 645311 0 FreeSans 320 0 0 0 gpio1_7_oe_n
port 984 nsew signal input
flabel metal3 s 677000 647022 677300 647142 0 FreeSans 320 0 0 0 gpio1_7_tie_lo_esd
port 985 nsew signal output
flabel metal3 s 677000 648625 677300 648691 0 FreeSans 320 0 0 0 gpio1_7_inp_dis
port 986 nsew signal input
flabel metal3 s 677000 650957 677300 651031 0 FreeSans 320 0 0 0 gpio1_7_enable_vddio
port 987 nsew signal input
flabel metal3 s 677000 652601 677300 652667 0 FreeSans 320 0 0 0 gpio1_7_vtrip_sel
port 988 nsew signal input
flabel metal3 s 677000 656747 677300 656813 0 FreeSans 320 0 0 0 gpio1_7_ib_mode_sel[1]
port 989 nsew signal input
flabel metal3 s 677000 652771 677300 652837 0 FreeSans 320 0 0 0 gpio1_7_ib_mode_sel[0]
port 990 nsew signal input
flabel metal3 s 677000 655309 677300 655375 0 FreeSans 320 0 0 0 gpio1_7_out
port 991 nsew signal input
flabel metal3 s 677000 660893 677300 660959 0 FreeSans 320 0 0 0 gpio1_7_slew_ctl[1]
port 992 nsew signal input
flabel metal3 s 677000 656917 677300 656983 0 FreeSans 320 0 0 0 gpio1_7_slew_ctl[0]
port 993 nsew signal input
flabel metal3 s 677000 657087 677300 657153 0 FreeSans 320 0 0 0 gpio1_7_analog_pol
port 994 nsew signal input
flabel metal3 s 677000 659803 677300 659869 0 FreeSans 320 0 0 0 gpio1_7_analog_sel
port 995 nsew signal input
flabel metal3 s 677000 661063 677300 661129 0 FreeSans 320 0 0 0 gpio1_7_hys_trim
port 996 nsew signal input
flabel metal3 s 677000 661327 677300 661393 0 FreeSans 320 0 0 0 gpio1_7_vinref
port 997 nsew signal input
flabel metal3 s 677000 664663 677300 664729 0 FreeSans 320 0 0 0 gpio1_7_hld_ovr
port 998 nsew signal input
flabel metal3 s 677000 665258 677300 665324 0 FreeSans 320 0 0 0 gpio1_7_in_h
port 999 nsew signal output
flabel metal3 s 677000 665707 677300 665773 0 FreeSans 320 0 0 0 gpio1_7_enable_h
port 1000 nsew signal input
flabel metal3 s 677000 666058 677300 666124 0 FreeSans 320 0 0 0 gpio1_7_in
port 1001 nsew signal output
flabel metal3 s 677000 666207 677300 666273 0 FreeSans 320 0 0 0 gpio1_7_hld_h_n
port 1002 nsew signal input
flabel metal3 s 677000 668380 677300 668446 0 FreeSans 320 0 0 0 gpio1_7_enable_vdda_h
port 1003 nsew signal input
flabel metal3 s 677000 668511 677300 668577 0 FreeSans 320 0 0 0 gpio1_7_analog_en
port 1004 nsew signal input
flabel metal3 s 677000 668712 677300 668778 0 FreeSans 320 0 0 0 gpio1_7_enable_inp_h
port 1005 nsew signal input
flabel metal3 s 677000 668927 677300 669047 0 FreeSans 320 0 0 0 gpio1_7_enable_vswitch_h
port 1006 nsew signal input
flabel metal3 s 677000 669503 677300 669623 0 FreeSans 320 0 0 0 gpio1_7_pad_a_noesd_h
port 1007 nsew signal bidirectional
flabel metal3 s 677000 669760 677300 669879 0 FreeSans 320 0 0 0 gpio1_7_pad_a_esd_0_h
port 1008 nsew signal bidirectional
flabel metal3 s 677000 670014 677300 670134 0 FreeSans 320 0 0 0 gpio1_7_pad_a_esd_1_h
port 1009 nsew signal bidirectional
flabel metal3 s 677000 640328 677300 640398 0 FreeSans 320 0 0 0 gpio1_7_zero
port 1010 nsew signal output
flabel metal3 s 677000 639878 677300 639948 0 FreeSans 320 0 0 0 gpio1_7_one
port 1011 nsew signal output
flabel metal3 s 676758 758528 677058 758598 0 FreeSans 320 0 0 0 gpio2_0_tie_lo_esd
port 1012 nsew signal output
flabel metal3 s 676762 759106 677062 759176 0 FreeSans 320 0 0 0 gpio2_0_in
port 1013 nsew signal output
flabel metal3 s 676758 758826 677058 758896 0 FreeSans 320 0 0 0 gpio2_0_tie_hi_esd
port 1014 nsew signal output
flabel metal3 s 676758 759418 677058 759488 0 FreeSans 320 0 0 0 gpio2_0_enable_vddio
port 1015 nsew signal input
flabel metal3 s 676758 759692 677058 759762 0 FreeSans 320 0 0 0 gpio2_0_slow
port 1016 nsew signal input
flabel metal3 s 676758 759982 677058 760110 0 FreeSans 320 0 0 0 gpio2_0_pad_a_esd_0_h
port 1017 nsew signal bidirectional
flabel metal3 s 676758 761412 677058 761542 0 FreeSans 320 0 0 0 gpio2_0_pad_a_esd_1_h
port 1018 nsew signal bidirectional
flabel metal3 s 676758 762422 677058 762636 0 FreeSans 320 0 0 0 gpio2_0_pad_a_noesd_h
port 1019 nsew signal bidirectional
flabel metal3 s 676758 763198 677058 763268 0 FreeSans 320 0 0 0 gpio2_0_analog_en
port 1020 nsew signal input
flabel metal3 s 676758 765958 677058 766028 0 FreeSans 320 0 0 0 gpio2_0_analog_pol
port 1021 nsew signal input
flabel metal3 s 676758 766538 677058 766608 0 FreeSans 320 0 0 0 gpio2_0_inp_dis
port 1022 nsew signal input
flabel metal3 s 676758 767704 677058 767774 0 FreeSans 320 0 0 0 gpio2_0_enable_inp_h
port 1023 nsew signal input
flabel metal3 s 676758 768160 677058 768230 0 FreeSans 320 0 0 0 gpio2_0_enable_h
port 1024 nsew signal input
flabel metal3 s 676758 768614 677058 768684 0 FreeSans 320 0 0 0 gpio2_0_hld_h_n
port 1025 nsew signal input
flabel metal3 s 676758 769232 677058 769302 0 FreeSans 320 0 0 0 gpio2_0_analog_sel
port 1026 nsew signal input
flabel metal3 s 676758 769676 677058 769746 0 FreeSans 320 0 0 0 gpio2_0_dm[2]
port 1027 nsew signal input
flabel metal3 s 676758 762002 677058 762072 0 FreeSans 320 0 0 0 gpio2_0_dm[1]
port 1028 nsew signal input
flabel metal3 s 676758 765410 677058 765480 0 FreeSans 320 0 0 0 gpio2_0_dm[0]
port 1029 nsew signal input
flabel metal3 s 676758 770160 677058 770230 0 FreeSans 320 0 0 0 gpio2_0_hld_ovr
port 1030 nsew signal input
flabel metal3 s 676758 770932 677058 771002 0 FreeSans 320 0 0 0 gpio2_0_out
port 1031 nsew signal input
flabel metal3 s 676758 772132 677058 772202 0 FreeSans 320 0 0 0 gpio2_0_enable_vswitch_h
port 1032 nsew signal input
flabel metal3 s 676758 772852 677058 772922 0 FreeSans 320 0 0 0 gpio2_0_enable_vdda_h
port 1033 nsew signal input
flabel metal3 s 676758 773714 677058 773784 0 FreeSans 320 0 0 0 gpio2_0_vtrip_sel
port 1034 nsew signal input
flabel metal3 s 676758 774058 677058 774128 0 FreeSans 320 0 0 0 gpio2_0_ib_mode_sel
port 1035 nsew signal input
flabel metal3 s 676758 774468 677058 774538 0 FreeSans 320 0 0 0 gpio2_0_oe_n
port 1036 nsew signal input
flabel metal3 s 676758 774996 677058 775120 0 FreeSans 320 0 0 0 gpio2_0_in_h
port 1037 nsew signal output
flabel metal3 s 676758 757328 677058 757398 0 FreeSans 320 0 0 0 gpio2_0_zero
port 1038 nsew signal output
flabel metal3 s 676758 756878 677058 756948 0 FreeSans 320 0 0 0 gpio2_0_one
port 1039 nsew signal output
flabel metal3 s 676758 779528 677058 779598 0 FreeSans 320 0 0 0 gpio2_1_tie_lo_esd
port 1040 nsew signal output
flabel metal3 s 676762 780106 677062 780176 0 FreeSans 320 0 0 0 gpio2_1_in
port 1041 nsew signal output
flabel metal3 s 676758 779826 677058 779896 0 FreeSans 320 0 0 0 gpio2_1_tie_hi_esd
port 1042 nsew signal output
flabel metal3 s 676758 780418 677058 780488 0 FreeSans 320 0 0 0 gpio2_1_enable_vddio
port 1043 nsew signal input
flabel metal3 s 676758 780692 677058 780762 0 FreeSans 320 0 0 0 gpio2_1_slow
port 1044 nsew signal input
flabel metal3 s 676758 780982 677058 781110 0 FreeSans 320 0 0 0 gpio2_1_pad_a_esd_0_h
port 1045 nsew signal bidirectional
flabel metal3 s 676758 782412 677058 782542 0 FreeSans 320 0 0 0 gpio2_1_pad_a_esd_1_h
port 1046 nsew signal bidirectional
flabel metal3 s 676758 783422 677058 783636 0 FreeSans 320 0 0 0 gpio2_1_pad_a_noesd_h
port 1047 nsew signal bidirectional
flabel metal3 s 676758 784198 677058 784268 0 FreeSans 320 0 0 0 gpio2_1_analog_en
port 1048 nsew signal input
flabel metal3 s 676758 786958 677058 787028 0 FreeSans 320 0 0 0 gpio2_1_analog_pol
port 1049 nsew signal input
flabel metal3 s 676758 787538 677058 787608 0 FreeSans 320 0 0 0 gpio2_1_inp_dis
port 1050 nsew signal input
flabel metal3 s 676758 788704 677058 788774 0 FreeSans 320 0 0 0 gpio2_1_enable_inp_h
port 1051 nsew signal input
flabel metal3 s 676758 789160 677058 789230 0 FreeSans 320 0 0 0 gpio2_1_enable_h
port 1052 nsew signal input
flabel metal3 s 676758 789614 677058 789684 0 FreeSans 320 0 0 0 gpio2_1_hld_h_n
port 1053 nsew signal input
flabel metal3 s 676758 790232 677058 790302 0 FreeSans 320 0 0 0 gpio2_1_analog_sel
port 1054 nsew signal input
flabel metal3 s 676758 790676 677058 790746 0 FreeSans 320 0 0 0 gpio2_1_dm[2]
port 1055 nsew signal input
flabel metal3 s 676758 783002 677058 783072 0 FreeSans 320 0 0 0 gpio2_1_dm[1]
port 1056 nsew signal input
flabel metal3 s 676758 786410 677058 786480 0 FreeSans 320 0 0 0 gpio2_1_dm[0]
port 1057 nsew signal input
flabel metal3 s 676758 791160 677058 791230 0 FreeSans 320 0 0 0 gpio2_1_hld_ovr
port 1058 nsew signal input
flabel metal3 s 676758 791932 677058 792002 0 FreeSans 320 0 0 0 gpio2_1_out
port 1059 nsew signal input
flabel metal3 s 676758 793132 677058 793202 0 FreeSans 320 0 0 0 gpio2_1_enable_vswitch_h
port 1060 nsew signal input
flabel metal3 s 676758 793852 677058 793922 0 FreeSans 320 0 0 0 gpio2_1_enable_vdda_h
port 1061 nsew signal input
flabel metal3 s 676758 794714 677058 794784 0 FreeSans 320 0 0 0 gpio2_1_vtrip_sel
port 1062 nsew signal input
flabel metal3 s 676758 795058 677058 795128 0 FreeSans 320 0 0 0 gpio2_1_ib_mode_sel
port 1063 nsew signal input
flabel metal3 s 676758 795468 677058 795538 0 FreeSans 320 0 0 0 gpio2_1_oe_n
port 1064 nsew signal input
flabel metal3 s 676758 795996 677058 796120 0 FreeSans 320 0 0 0 gpio2_1_in_h
port 1065 nsew signal output
flabel metal3 s 676758 778328 677058 778398 0 FreeSans 320 0 0 0 gpio2_1_zero
port 1066 nsew signal output
flabel metal3 s 676758 777878 677058 777948 0 FreeSans 320 0 0 0 gpio2_1_one
port 1067 nsew signal output
flabel metal3 s 676758 800528 677058 800598 0 FreeSans 320 0 0 0 gpio2_2_tie_lo_esd
port 1068 nsew signal output
flabel metal3 s 676762 801106 677062 801176 0 FreeSans 320 0 0 0 gpio2_2_in
port 1069 nsew signal output
flabel metal3 s 676758 800826 677058 800896 0 FreeSans 320 0 0 0 gpio2_2_tie_hi_esd
port 1070 nsew signal output
flabel metal3 s 676758 801418 677058 801488 0 FreeSans 320 0 0 0 gpio2_2_enable_vddio
port 1071 nsew signal input
flabel metal3 s 676758 801692 677058 801762 0 FreeSans 320 0 0 0 gpio2_2_slow
port 1072 nsew signal input
flabel metal3 s 676758 801982 677058 802110 0 FreeSans 320 0 0 0 gpio2_2_pad_a_esd_0_h
port 1073 nsew signal bidirectional
flabel metal3 s 676758 803412 677058 803542 0 FreeSans 320 0 0 0 gpio2_2_pad_a_esd_1_h
port 1074 nsew signal bidirectional
flabel metal3 s 676758 804422 677058 804636 0 FreeSans 320 0 0 0 gpio2_2_pad_a_noesd_h
port 1075 nsew signal bidirectional
flabel metal3 s 676758 805198 677058 805268 0 FreeSans 320 0 0 0 gpio2_2_analog_en
port 1076 nsew signal input
flabel metal3 s 676758 807958 677058 808028 0 FreeSans 320 0 0 0 gpio2_2_analog_pol
port 1077 nsew signal input
flabel metal3 s 676758 808538 677058 808608 0 FreeSans 320 0 0 0 gpio2_2_inp_dis
port 1078 nsew signal input
flabel metal3 s 676758 809704 677058 809774 0 FreeSans 320 0 0 0 gpio2_2_enable_inp_h
port 1079 nsew signal input
flabel metal3 s 676758 810160 677058 810230 0 FreeSans 320 0 0 0 gpio2_2_enable_h
port 1080 nsew signal input
flabel metal3 s 676758 810614 677058 810684 0 FreeSans 320 0 0 0 gpio2_2_hld_h_n
port 1081 nsew signal input
flabel metal3 s 676758 811232 677058 811302 0 FreeSans 320 0 0 0 gpio2_2_analog_sel
port 1082 nsew signal input
flabel metal3 s 676758 811676 677058 811746 0 FreeSans 320 0 0 0 gpio2_2_dm[2]
port 1083 nsew signal input
flabel metal3 s 676758 804002 677058 804072 0 FreeSans 320 0 0 0 gpio2_2_dm[1]
port 1084 nsew signal input
flabel metal3 s 676758 807410 677058 807480 0 FreeSans 320 0 0 0 gpio2_2_dm[0]
port 1085 nsew signal input
flabel metal3 s 676758 812160 677058 812230 0 FreeSans 320 0 0 0 gpio2_2_hld_ovr
port 1086 nsew signal input
flabel metal3 s 676758 812932 677058 813002 0 FreeSans 320 0 0 0 gpio2_2_out
port 1087 nsew signal input
flabel metal3 s 676758 814132 677058 814202 0 FreeSans 320 0 0 0 gpio2_2_enable_vswitch_h
port 1088 nsew signal input
flabel metal3 s 676758 814852 677058 814922 0 FreeSans 320 0 0 0 gpio2_2_enable_vdda_h
port 1089 nsew signal input
flabel metal3 s 676758 815714 677058 815784 0 FreeSans 320 0 0 0 gpio2_2_vtrip_sel
port 1090 nsew signal input
flabel metal3 s 676758 816058 677058 816128 0 FreeSans 320 0 0 0 gpio2_2_ib_mode_sel
port 1091 nsew signal input
flabel metal3 s 676758 816468 677058 816538 0 FreeSans 320 0 0 0 gpio2_2_oe_n
port 1092 nsew signal input
flabel metal3 s 676758 816996 677058 817120 0 FreeSans 320 0 0 0 gpio2_2_in_h
port 1093 nsew signal output
flabel metal3 s 676758 799328 677058 799398 0 FreeSans 320 0 0 0 gpio2_2_zero
port 1094 nsew signal output
flabel metal3 s 676758 798878 677058 798948 0 FreeSans 320 0 0 0 gpio2_2_one
port 1095 nsew signal output
flabel metal3 s 676758 821528 677058 821598 0 FreeSans 320 0 0 0 gpio2_3_tie_lo_esd
port 1096 nsew signal output
flabel metal3 s 676762 822106 677062 822176 0 FreeSans 320 0 0 0 gpio2_3_in
port 1097 nsew signal output
flabel metal3 s 676758 821826 677058 821896 0 FreeSans 320 0 0 0 gpio2_3_tie_hi_esd
port 1098 nsew signal output
flabel metal3 s 676758 822418 677058 822488 0 FreeSans 320 0 0 0 gpio2_3_enable_vddio
port 1099 nsew signal input
flabel metal3 s 676758 822692 677058 822762 0 FreeSans 320 0 0 0 gpio2_3_slow
port 1100 nsew signal input
flabel metal3 s 676758 822982 677058 823110 0 FreeSans 320 0 0 0 gpio2_3_pad_a_esd_0_h
port 1101 nsew signal bidirectional
flabel metal3 s 676758 824412 677058 824542 0 FreeSans 320 0 0 0 gpio2_3_pad_a_esd_1_h
port 1102 nsew signal bidirectional
flabel metal3 s 676758 825422 677058 825636 0 FreeSans 320 0 0 0 gpio2_3_pad_a_noesd_h
port 1103 nsew signal bidirectional
flabel metal3 s 676758 826198 677058 826268 0 FreeSans 320 0 0 0 gpio2_3_analog_en
port 1104 nsew signal input
flabel metal3 s 676758 828958 677058 829028 0 FreeSans 320 0 0 0 gpio2_3_analog_pol
port 1105 nsew signal input
flabel metal3 s 676758 829538 677058 829608 0 FreeSans 320 0 0 0 gpio2_3_inp_dis
port 1106 nsew signal input
flabel metal3 s 676758 830704 677058 830774 0 FreeSans 320 0 0 0 gpio2_3_enable_inp_h
port 1107 nsew signal input
flabel metal3 s 676758 831160 677058 831230 0 FreeSans 320 0 0 0 gpio2_3_enable_h
port 1108 nsew signal input
flabel metal3 s 676758 831614 677058 831684 0 FreeSans 320 0 0 0 gpio2_3_hld_h_n
port 1109 nsew signal input
flabel metal3 s 676758 832232 677058 832302 0 FreeSans 320 0 0 0 gpio2_3_analog_sel
port 1110 nsew signal input
flabel metal3 s 676758 832676 677058 832746 0 FreeSans 320 0 0 0 gpio2_3_dm[2]
port 1111 nsew signal input
flabel metal3 s 676758 825002 677058 825072 0 FreeSans 320 0 0 0 gpio2_3_dm[1]
port 1112 nsew signal input
flabel metal3 s 676758 828410 677058 828480 0 FreeSans 320 0 0 0 gpio2_3_dm[0]
port 1113 nsew signal input
flabel metal3 s 676758 833160 677058 833230 0 FreeSans 320 0 0 0 gpio2_3_hld_ovr
port 1114 nsew signal input
flabel metal3 s 676758 833932 677058 834002 0 FreeSans 320 0 0 0 gpio2_3_out
port 1115 nsew signal input
flabel metal3 s 676758 835132 677058 835202 0 FreeSans 320 0 0 0 gpio2_3_enable_vswitch_h
port 1116 nsew signal input
flabel metal3 s 676758 835852 677058 835922 0 FreeSans 320 0 0 0 gpio2_3_enable_vdda_h
port 1117 nsew signal input
flabel metal3 s 676758 836714 677058 836784 0 FreeSans 320 0 0 0 gpio2_3_vtrip_sel
port 1118 nsew signal input
flabel metal3 s 676758 837058 677058 837128 0 FreeSans 320 0 0 0 gpio2_3_ib_mode_sel
port 1119 nsew signal input
flabel metal3 s 676758 837468 677058 837538 0 FreeSans 320 0 0 0 gpio2_3_oe_n
port 1120 nsew signal input
flabel metal3 s 676758 837996 677058 838120 0 FreeSans 320 0 0 0 gpio2_3_in_h
port 1121 nsew signal output
flabel metal3 s 676758 820328 677058 820398 0 FreeSans 320 0 0 0 gpio2_3_zero
port 1122 nsew signal output
flabel metal3 s 676758 819878 677058 819948 0 FreeSans 320 0 0 0 gpio2_3_one
port 1123 nsew signal output
flabel metal3 s 676758 862528 677058 862598 0 FreeSans 320 0 0 0 gpio2_4_tie_lo_esd
port 1124 nsew signal output
flabel metal3 s 676762 863106 677062 863176 0 FreeSans 320 0 0 0 gpio2_4_in
port 1125 nsew signal output
flabel metal3 s 676758 862826 677058 862896 0 FreeSans 320 0 0 0 gpio2_4_tie_hi_esd
port 1126 nsew signal output
flabel metal3 s 676758 863418 677058 863488 0 FreeSans 320 0 0 0 gpio2_4_enable_vddio
port 1127 nsew signal input
flabel metal3 s 676758 863692 677058 863762 0 FreeSans 320 0 0 0 gpio2_4_slow
port 1128 nsew signal input
flabel metal3 s 676758 863982 677058 864110 0 FreeSans 320 0 0 0 gpio2_4_pad_a_esd_0_h
port 1129 nsew signal bidirectional
flabel metal3 s 676758 865412 677058 865542 0 FreeSans 320 0 0 0 gpio2_4_pad_a_esd_1_h
port 1130 nsew signal bidirectional
flabel metal3 s 676758 866422 677058 866636 0 FreeSans 320 0 0 0 gpio2_4_pad_a_noesd_h
port 1131 nsew signal bidirectional
flabel metal3 s 676758 867198 677058 867268 0 FreeSans 320 0 0 0 gpio2_4_analog_en
port 1132 nsew signal input
flabel metal3 s 676758 869958 677058 870028 0 FreeSans 320 0 0 0 gpio2_4_analog_pol
port 1133 nsew signal input
flabel metal3 s 676758 870538 677058 870608 0 FreeSans 320 0 0 0 gpio2_4_inp_dis
port 1134 nsew signal input
flabel metal3 s 676758 871704 677058 871774 0 FreeSans 320 0 0 0 gpio2_4_enable_inp_h
port 1135 nsew signal input
flabel metal3 s 676758 872160 677058 872230 0 FreeSans 320 0 0 0 gpio2_4_enable_h
port 1136 nsew signal input
flabel metal3 s 676758 872614 677058 872684 0 FreeSans 320 0 0 0 gpio2_4_hld_h_n
port 1137 nsew signal input
flabel metal3 s 676758 873232 677058 873302 0 FreeSans 320 0 0 0 gpio2_4_analog_sel
port 1138 nsew signal input
flabel metal3 s 676758 873676 677058 873746 0 FreeSans 320 0 0 0 gpio2_4_dm[2]
port 1139 nsew signal input
flabel metal3 s 676758 866002 677058 866072 0 FreeSans 320 0 0 0 gpio2_4_dm[1]
port 1140 nsew signal input
flabel metal3 s 676758 869410 677058 869480 0 FreeSans 320 0 0 0 gpio2_4_dm[0]
port 1141 nsew signal input
flabel metal3 s 676758 874160 677058 874230 0 FreeSans 320 0 0 0 gpio2_4_hld_ovr
port 1142 nsew signal input
flabel metal3 s 676758 874932 677058 875002 0 FreeSans 320 0 0 0 gpio2_4_out
port 1143 nsew signal input
flabel metal3 s 676758 876132 677058 876202 0 FreeSans 320 0 0 0 gpio2_4_enable_vswitch_h
port 1144 nsew signal input
flabel metal3 s 676758 876852 677058 876922 0 FreeSans 320 0 0 0 gpio2_4_enable_vdda_h
port 1145 nsew signal input
flabel metal3 s 676758 877714 677058 877784 0 FreeSans 320 0 0 0 gpio2_4_vtrip_sel
port 1146 nsew signal input
flabel metal3 s 676758 878058 677058 878128 0 FreeSans 320 0 0 0 gpio2_4_ib_mode_sel
port 1147 nsew signal input
flabel metal3 s 676758 878468 677058 878538 0 FreeSans 320 0 0 0 gpio2_4_oe_n
port 1148 nsew signal input
flabel metal3 s 676758 878996 677058 879120 0 FreeSans 320 0 0 0 gpio2_4_in_h
port 1149 nsew signal output
flabel metal3 s 676758 861328 677058 861398 0 FreeSans 320 0 0 0 gpio2_4_zero
port 1150 nsew signal output
flabel metal3 s 676758 860878 677058 860948 0 FreeSans 320 0 0 0 gpio2_4_one
port 1151 nsew signal output
flabel metal3 s 676758 883528 677058 883598 0 FreeSans 320 0 0 0 gpio2_5_tie_lo_esd
port 1152 nsew signal output
flabel metal3 s 676762 884106 677062 884176 0 FreeSans 320 0 0 0 gpio2_5_in
port 1153 nsew signal output
flabel metal3 s 676758 883826 677058 883896 0 FreeSans 320 0 0 0 gpio2_5_tie_hi_esd
port 1154 nsew signal output
flabel metal3 s 676758 884418 677058 884488 0 FreeSans 320 0 0 0 gpio2_5_enable_vddio
port 1155 nsew signal input
flabel metal3 s 676758 884692 677058 884762 0 FreeSans 320 0 0 0 gpio2_5_slow
port 1156 nsew signal input
flabel metal3 s 676758 884982 677058 885110 0 FreeSans 320 0 0 0 gpio2_5_pad_a_esd_0_h
port 1157 nsew signal bidirectional
flabel metal3 s 676758 886412 677058 886542 0 FreeSans 320 0 0 0 gpio2_5_pad_a_esd_1_h
port 1158 nsew signal bidirectional
flabel metal3 s 676758 887422 677058 887636 0 FreeSans 320 0 0 0 gpio2_5_pad_a_noesd_h
port 1159 nsew signal bidirectional
flabel metal3 s 676758 888198 677058 888268 0 FreeSans 320 0 0 0 gpio2_5_analog_en
port 1160 nsew signal input
flabel metal3 s 676758 890958 677058 891028 0 FreeSans 320 0 0 0 gpio2_5_analog_pol
port 1161 nsew signal input
flabel metal3 s 676758 891538 677058 891608 0 FreeSans 320 0 0 0 gpio2_5_inp_dis
port 1162 nsew signal input
flabel metal3 s 676758 892704 677058 892774 0 FreeSans 320 0 0 0 gpio2_5_enable_inp_h
port 1163 nsew signal input
flabel metal3 s 676758 893160 677058 893230 0 FreeSans 320 0 0 0 gpio2_5_enable_h
port 1164 nsew signal input
flabel metal3 s 676758 893614 677058 893684 0 FreeSans 320 0 0 0 gpio2_5_hld_h_n
port 1165 nsew signal input
flabel metal3 s 676758 894232 677058 894302 0 FreeSans 320 0 0 0 gpio2_5_analog_sel
port 1166 nsew signal input
flabel metal3 s 676758 894676 677058 894746 0 FreeSans 320 0 0 0 gpio2_5_dm[2]
port 1167 nsew signal input
flabel metal3 s 676758 887002 677058 887072 0 FreeSans 320 0 0 0 gpio2_5_dm[1]
port 1168 nsew signal input
flabel metal3 s 676758 890410 677058 890480 0 FreeSans 320 0 0 0 gpio2_5_dm[0]
port 1169 nsew signal input
flabel metal3 s 676758 895160 677058 895230 0 FreeSans 320 0 0 0 gpio2_5_hld_ovr
port 1170 nsew signal input
flabel metal3 s 676758 895932 677058 896002 0 FreeSans 320 0 0 0 gpio2_5_out
port 1171 nsew signal input
flabel metal3 s 676758 897132 677058 897202 0 FreeSans 320 0 0 0 gpio2_5_enable_vswitch_h
port 1172 nsew signal input
flabel metal3 s 676758 897852 677058 897922 0 FreeSans 320 0 0 0 gpio2_5_enable_vdda_h
port 1173 nsew signal input
flabel metal3 s 676758 898714 677058 898784 0 FreeSans 320 0 0 0 gpio2_5_vtrip_sel
port 1174 nsew signal input
flabel metal3 s 676758 899058 677058 899128 0 FreeSans 320 0 0 0 gpio2_5_ib_mode_sel
port 1175 nsew signal input
flabel metal3 s 676758 899468 677058 899538 0 FreeSans 320 0 0 0 gpio2_5_oe_n
port 1176 nsew signal input
flabel metal3 s 676758 899996 677058 900120 0 FreeSans 320 0 0 0 gpio2_5_in_h
port 1177 nsew signal output
flabel metal3 s 676758 882328 677058 882398 0 FreeSans 320 0 0 0 gpio2_5_zero
port 1178 nsew signal output
flabel metal3 s 676758 881878 677058 881948 0 FreeSans 320 0 0 0 gpio2_5_one
port 1179 nsew signal output
flabel metal3 s 676758 904528 677058 904598 0 FreeSans 320 0 0 0 gpio2_6_tie_lo_esd
port 1180 nsew signal output
flabel metal3 s 676762 905106 677062 905176 0 FreeSans 320 0 0 0 gpio2_6_in
port 1181 nsew signal output
flabel metal3 s 676758 904826 677058 904896 0 FreeSans 320 0 0 0 gpio2_6_tie_hi_esd
port 1182 nsew signal output
flabel metal3 s 676758 905418 677058 905488 0 FreeSans 320 0 0 0 gpio2_6_enable_vddio
port 1183 nsew signal input
flabel metal3 s 676758 905692 677058 905762 0 FreeSans 320 0 0 0 gpio2_6_slow
port 1184 nsew signal input
flabel metal3 s 676758 905982 677058 906110 0 FreeSans 320 0 0 0 gpio2_6_pad_a_esd_0_h
port 1185 nsew signal bidirectional
flabel metal3 s 676758 907412 677058 907542 0 FreeSans 320 0 0 0 gpio2_6_pad_a_esd_1_h
port 1186 nsew signal bidirectional
flabel metal3 s 676758 908422 677058 908636 0 FreeSans 320 0 0 0 gpio2_6_pad_a_noesd_h
port 1187 nsew signal bidirectional
flabel metal3 s 676758 909198 677058 909268 0 FreeSans 320 0 0 0 gpio2_6_analog_en
port 1188 nsew signal input
flabel metal3 s 676758 911958 677058 912028 0 FreeSans 320 0 0 0 gpio2_6_analog_pol
port 1189 nsew signal input
flabel metal3 s 676758 912538 677058 912608 0 FreeSans 320 0 0 0 gpio2_6_inp_dis
port 1190 nsew signal input
flabel metal3 s 676758 913704 677058 913774 0 FreeSans 320 0 0 0 gpio2_6_enable_inp_h
port 1191 nsew signal input
flabel metal3 s 676758 914160 677058 914230 0 FreeSans 320 0 0 0 gpio2_6_enable_h
port 1192 nsew signal input
flabel metal3 s 676758 914614 677058 914684 0 FreeSans 320 0 0 0 gpio2_6_hld_h_n
port 1193 nsew signal input
flabel metal3 s 676758 915232 677058 915302 0 FreeSans 320 0 0 0 gpio2_6_analog_sel
port 1194 nsew signal input
flabel metal3 s 676758 915676 677058 915746 0 FreeSans 320 0 0 0 gpio2_6_dm[2]
port 1195 nsew signal input
flabel metal3 s 676758 908002 677058 908072 0 FreeSans 320 0 0 0 gpio2_6_dm[1]
port 1196 nsew signal input
flabel metal3 s 676758 911410 677058 911480 0 FreeSans 320 0 0 0 gpio2_6_dm[0]
port 1197 nsew signal input
flabel metal3 s 676758 916160 677058 916230 0 FreeSans 320 0 0 0 gpio2_6_hld_ovr
port 1198 nsew signal input
flabel metal3 s 676758 916932 677058 917002 0 FreeSans 320 0 0 0 gpio2_6_out
port 1199 nsew signal input
flabel metal3 s 676758 918132 677058 918202 0 FreeSans 320 0 0 0 gpio2_6_enable_vswitch_h
port 1200 nsew signal input
flabel metal3 s 676758 918852 677058 918922 0 FreeSans 320 0 0 0 gpio2_6_enable_vdda_h
port 1201 nsew signal input
flabel metal3 s 676758 919714 677058 919784 0 FreeSans 320 0 0 0 gpio2_6_vtrip_sel
port 1202 nsew signal input
flabel metal3 s 676758 920058 677058 920128 0 FreeSans 320 0 0 0 gpio2_6_ib_mode_sel
port 1203 nsew signal input
flabel metal3 s 676758 920468 677058 920538 0 FreeSans 320 0 0 0 gpio2_6_oe_n
port 1204 nsew signal input
flabel metal3 s 676758 920996 677058 921120 0 FreeSans 320 0 0 0 gpio2_6_in_h
port 1205 nsew signal output
flabel metal3 s 676758 903328 677058 903398 0 FreeSans 320 0 0 0 gpio2_6_zero
port 1206 nsew signal output
flabel metal3 s 676758 902878 677058 902948 0 FreeSans 320 0 0 0 gpio2_6_one
port 1207 nsew signal output
flabel metal3 s 676758 925528 677058 925598 0 FreeSans 320 0 0 0 gpio2_7_tie_lo_esd
port 1208 nsew signal output
flabel metal3 s 676762 926106 677062 926176 0 FreeSans 320 0 0 0 gpio2_7_in
port 1209 nsew signal output
flabel metal3 s 676758 925826 677058 925896 0 FreeSans 320 0 0 0 gpio2_7_tie_hi_esd
port 1210 nsew signal output
flabel metal3 s 676758 926418 677058 926488 0 FreeSans 320 0 0 0 gpio2_7_enable_vddio
port 1211 nsew signal input
flabel metal3 s 676758 926692 677058 926762 0 FreeSans 320 0 0 0 gpio2_7_slow
port 1212 nsew signal input
flabel metal3 s 676758 926982 677058 927110 0 FreeSans 320 0 0 0 gpio2_7_pad_a_esd_0_h
port 1213 nsew signal bidirectional
flabel metal3 s 676758 928412 677058 928542 0 FreeSans 320 0 0 0 gpio2_7_pad_a_esd_1_h
port 1214 nsew signal bidirectional
flabel metal3 s 676758 929422 677058 929636 0 FreeSans 320 0 0 0 gpio2_7_pad_a_noesd_h
port 1215 nsew signal bidirectional
flabel metal3 s 676758 930198 677058 930268 0 FreeSans 320 0 0 0 gpio2_7_analog_en
port 1216 nsew signal input
flabel metal3 s 676758 932958 677058 933028 0 FreeSans 320 0 0 0 gpio2_7_analog_pol
port 1217 nsew signal input
flabel metal3 s 676758 933538 677058 933608 0 FreeSans 320 0 0 0 gpio2_7_inp_dis
port 1218 nsew signal input
flabel metal3 s 676758 934704 677058 934774 0 FreeSans 320 0 0 0 gpio2_7_enable_inp_h
port 1219 nsew signal input
flabel metal3 s 676758 935160 677058 935230 0 FreeSans 320 0 0 0 gpio2_7_enable_h
port 1220 nsew signal input
flabel metal3 s 676758 935614 677058 935684 0 FreeSans 320 0 0 0 gpio2_7_hld_h_n
port 1221 nsew signal input
flabel metal3 s 676758 936232 677058 936302 0 FreeSans 320 0 0 0 gpio2_7_analog_sel
port 1222 nsew signal input
flabel metal3 s 676758 936676 677058 936746 0 FreeSans 320 0 0 0 gpio2_7_dm[2]
port 1223 nsew signal input
flabel metal3 s 676758 929002 677058 929072 0 FreeSans 320 0 0 0 gpio2_7_dm[1]
port 1224 nsew signal input
flabel metal3 s 676758 932410 677058 932480 0 FreeSans 320 0 0 0 gpio2_7_dm[0]
port 1225 nsew signal input
flabel metal3 s 676758 937160 677058 937230 0 FreeSans 320 0 0 0 gpio2_7_hld_ovr
port 1226 nsew signal input
flabel metal3 s 676758 937932 677058 938002 0 FreeSans 320 0 0 0 gpio2_7_out
port 1227 nsew signal input
flabel metal3 s 676758 939132 677058 939202 0 FreeSans 320 0 0 0 gpio2_7_enable_vswitch_h
port 1228 nsew signal input
flabel metal3 s 676758 939852 677058 939922 0 FreeSans 320 0 0 0 gpio2_7_enable_vdda_h
port 1229 nsew signal input
flabel metal3 s 676758 940714 677058 940784 0 FreeSans 320 0 0 0 gpio2_7_vtrip_sel
port 1230 nsew signal input
flabel metal3 s 676758 941058 677058 941128 0 FreeSans 320 0 0 0 gpio2_7_ib_mode_sel
port 1231 nsew signal input
flabel metal3 s 676758 941468 677058 941538 0 FreeSans 320 0 0 0 gpio2_7_oe_n
port 1232 nsew signal input
flabel metal3 s 676758 941996 677058 942120 0 FreeSans 320 0 0 0 gpio2_7_in_h
port 1233 nsew signal output
flabel metal3 s 676758 924328 677058 924398 0 FreeSans 320 0 0 0 gpio2_7_zero
port 1234 nsew signal output
flabel metal3 s 676758 923878 677058 923948 0 FreeSans 320 0 0 0 gpio2_7_one
port 1235 nsew signal output
flabel metal3 s 676700 989586 677000 989646 0 FreeSans 320 0 0 0 muxsplit_ne_hld_vdda_h_n
port 1236 nsew signal input
flabel metal3 s 676700 990466 677000 990526 0 FreeSans 320 0 0 0 muxsplit_ne_enable_vdda_h
port 1237 nsew signal input
flabel metal3 s 676700 994088 677000 994148 0 FreeSans 320 0 0 0 muxsplit_ne_switch_aa_sl
port 1238 nsew signal input
flabel metal3 s 676700 994340 677000 994400 0 FreeSans 320 0 0 0 muxsplit_ne_switch_aa_s0
port 1239 nsew signal input
flabel metal3 s 676700 994592 677000 994652 0 FreeSans 320 0 0 0 muxsplit_ne_switch_bb_s0
port 1240 nsew signal input
flabel metal3 s 676700 994844 677000 994904 0 FreeSans 320 0 0 0 muxsplit_ne_switch_bb_sl
port 1241 nsew signal input
flabel metal3 s 676700 995096 677000 995156 0 FreeSans 320 0 0 0 muxsplit_ne_switch_bb_sr
port 1242 nsew signal input
flabel metal3 s 676700 995432 677000 995492 0 FreeSans 320 0 0 0 muxsplit_ne_switch_aa_sr
port 1243 nsew signal input
flabel metal2 s 651290 996690 651342 996890 0 FreeSans 320 90 0 0 gpio3_0_tie_lo_esd
port 1244 nsew signal output
flabel metal2 s 650990 996690 651042 996890 0 FreeSans 320 90 0 0 gpio3_0_in
port 1245 nsew signal output
flabel metal2 s 650688 996690 650740 996890 0 FreeSans 320 90 0 0 gpio3_0_tie_hi_esd
port 1246 nsew signal output
flabel metal2 s 650390 996690 650442 996890 0 FreeSans 320 90 0 0 gpio3_0_enable_vddio
port 1247 nsew signal input
flabel metal2 s 650090 996690 650142 996890 0 FreeSans 320 90 0 0 gpio3_0_slow
port 1248 nsew signal input
flabel metal2 s 649714 996690 649842 996890 0 FreeSans 320 90 0 0 gpio3_0_pad_a_esd_0_h
port 1249 nsew signal bidirectional
flabel metal2 s 648454 996690 648584 996890 0 FreeSans 320 90 0 0 gpio3_0_pad_a_esd_1_h
port 1250 nsew signal bidirectional
flabel metal2 s 647362 996690 647576 996890 0 FreeSans 320 90 0 0 gpio3_0_pad_a_noesd_h
port 1251 nsew signal bidirectional
flabel metal2 s 647058 996690 647110 996890 0 FreeSans 320 90 0 0 gpio3_0_analog_en
port 1252 nsew signal input
flabel metal2 s 644144 996690 644196 996890 0 FreeSans 320 90 0 0 gpio3_0_analog_pol
port 1253 nsew signal input
flabel metal2 s 643848 996690 643900 996890 0 FreeSans 320 90 0 0 gpio3_0_inp_dis
port 1254 nsew signal input
flabel metal2 s 642473 996690 642529 996890 0 FreeSans 320 90 0 0 gpio3_0_enable_inp_h
port 1255 nsew signal input
flabel metal2 s 641891 996690 641943 996890 0 FreeSans 320 90 0 0 gpio3_0_enable_h
port 1256 nsew signal input
flabel metal2 s 641162 996690 641214 996890 0 FreeSans 320 90 0 0 gpio3_0_hld_h_n
port 1257 nsew signal input
flabel metal2 s 640848 996690 640900 996890 0 FreeSans 320 90 0 0 gpio3_0_analog_sel
port 1258 nsew signal input
flabel metal2 s 640497 996690 640549 996890 0 FreeSans 320 90 0 0 gpio3_0_dm[2]
port 1259 nsew signal input
flabel metal2 s 648166 996690 648218 996890 0 FreeSans 320 90 0 0 gpio3_0_dm[1]
port 1260 nsew signal input
flabel metal2 s 644770 996690 644822 996890 0 FreeSans 320 90 0 0 gpio3_0_dm[0]
port 1261 nsew signal input
flabel metal2 s 640119 996690 640171 996890 0 FreeSans 320 90 0 0 gpio3_0_hld_ovr
port 1262 nsew signal input
flabel metal2 s 639270 996690 639322 996890 0 FreeSans 320 90 0 0 gpio3_0_out
port 1263 nsew signal input
flabel metal2 s 638061 996690 638113 996890 0 FreeSans 320 90 0 0 gpio3_0_enable_vswitch_h
port 1264 nsew signal input
flabel metal2 s 637350 996690 637402 996890 0 FreeSans 320 90 0 0 gpio3_0_enable_vdda_h
port 1265 nsew signal input
flabel metal2 s 636102 996690 636154 996890 0 FreeSans 320 90 0 0 gpio3_0_vtrip_sel
port 1266 nsew signal input
flabel metal2 s 635782 996690 635834 996890 0 FreeSans 320 90 0 0 gpio3_0_ib_mode_sel
port 1267 nsew signal input
flabel metal2 s 635468 996690 635520 996890 0 FreeSans 320 90 0 0 gpio3_0_oe_n
port 1268 nsew signal input
flabel metal2 s 634878 996690 635002 996890 0 FreeSans 320 90 0 0 gpio3_0_in_h
port 1269 nsew signal input
flabel metal2 s 652254 996690 652306 996890 0 FreeSans 320 90 0 0 gpio3_0_zero
port 1270 nsew signal output
flabel metal2 s 652616 996690 652668 996890 0 FreeSans 320 90 0 0 gpio3_0_one
port 1271 nsew signal output
flabel metal2 s 627290 996690 627342 996890 0 FreeSans 320 90 0 0 gpio3_1_tie_lo_esd
port 1272 nsew signal output
flabel metal2 s 626990 996690 627042 996890 0 FreeSans 320 90 0 0 gpio3_1_in
port 1273 nsew signal output
flabel metal2 s 626688 996690 626740 996890 0 FreeSans 320 90 0 0 gpio3_1_tie_hi_esd
port 1274 nsew signal output
flabel metal2 s 626390 996690 626442 996890 0 FreeSans 320 90 0 0 gpio3_1_enable_vddio
port 1275 nsew signal input
flabel metal2 s 626090 996690 626142 996890 0 FreeSans 320 90 0 0 gpio3_1_slow
port 1276 nsew signal input
flabel metal2 s 625714 996690 625842 996890 0 FreeSans 320 90 0 0 gpio3_1_pad_a_esd_0_h
port 1277 nsew signal bidirectional
flabel metal2 s 624454 996690 624584 996890 0 FreeSans 320 90 0 0 gpio3_1_pad_a_esd_1_h
port 1278 nsew signal bidirectional
flabel metal2 s 623362 996690 623576 996890 0 FreeSans 320 90 0 0 gpio3_1_pad_a_noesd_h
port 1279 nsew signal bidirectional
flabel metal2 s 623058 996690 623110 996890 0 FreeSans 320 90 0 0 gpio3_1_analog_en
port 1280 nsew signal input
flabel metal2 s 620144 996690 620196 996890 0 FreeSans 320 90 0 0 gpio3_1_analog_pol
port 1281 nsew signal input
flabel metal2 s 619848 996690 619900 996890 0 FreeSans 320 90 0 0 gpio3_1_inp_dis
port 1282 nsew signal input
flabel metal2 s 618473 996690 618529 996890 0 FreeSans 320 90 0 0 gpio3_1_enable_inp_h
port 1283 nsew signal input
flabel metal2 s 617891 996690 617943 996890 0 FreeSans 320 90 0 0 gpio3_1_enable_h
port 1284 nsew signal input
flabel metal2 s 617162 996690 617214 996890 0 FreeSans 320 90 0 0 gpio3_1_hld_h_n
port 1285 nsew signal input
flabel metal2 s 616848 996690 616900 996890 0 FreeSans 320 90 0 0 gpio3_1_analog_sel
port 1286 nsew signal input
flabel metal2 s 616497 996690 616549 996890 0 FreeSans 320 90 0 0 gpio3_1_dm[2]
port 1287 nsew signal input
flabel metal2 s 624166 996690 624218 996890 0 FreeSans 320 90 0 0 gpio3_1_dm[1]
port 1288 nsew signal input
flabel metal2 s 620770 996690 620822 996890 0 FreeSans 320 90 0 0 gpio3_1_dm[0]
port 1289 nsew signal input
flabel metal2 s 616119 996690 616171 996890 0 FreeSans 320 90 0 0 gpio3_1_hld_ovr
port 1290 nsew signal input
flabel metal2 s 615270 996690 615322 996890 0 FreeSans 320 90 0 0 gpio3_1_out
port 1291 nsew signal input
flabel metal2 s 614061 996690 614113 996890 0 FreeSans 320 90 0 0 gpio3_1_enable_vswitch_h
port 1292 nsew signal input
flabel metal2 s 613350 996690 613402 996890 0 FreeSans 320 90 0 0 gpio3_1_enable_vdda_h
port 1293 nsew signal input
flabel metal2 s 612102 996690 612154 996890 0 FreeSans 320 90 0 0 gpio3_1_vtrip_sel
port 1294 nsew signal input
flabel metal2 s 611782 996690 611834 996890 0 FreeSans 320 90 0 0 gpio3_1_ib_mode_sel
port 1295 nsew signal input
flabel metal2 s 611468 996690 611520 996890 0 FreeSans 320 90 0 0 gpio3_1_oe_n
port 1296 nsew signal input
flabel metal2 s 610878 996690 611002 996890 0 FreeSans 320 90 0 0 gpio3_1_in_h
port 1297 nsew signal input
flabel metal2 s 628254 996690 628306 996890 0 FreeSans 320 90 0 0 gpio3_1_zero
port 1298 nsew signal output
flabel metal2 s 628616 996690 628668 996890 0 FreeSans 320 90 0 0 gpio3_1_one
port 1299 nsew signal output
flabel metal2 s 603290 996690 603342 996890 0 FreeSans 320 90 0 0 gpio3_2_tie_lo_esd
port 1300 nsew signal output
flabel metal2 s 602990 996690 603042 996890 0 FreeSans 320 90 0 0 gpio3_2_in
port 1301 nsew signal output
flabel metal2 s 602688 996690 602740 996890 0 FreeSans 320 90 0 0 gpio3_2_tie_hi_esd
port 1302 nsew signal output
flabel metal2 s 602390 996690 602442 996890 0 FreeSans 320 90 0 0 gpio3_2_enable_vddio
port 1303 nsew signal input
flabel metal2 s 602090 996690 602142 996890 0 FreeSans 320 90 0 0 gpio3_2_slow
port 1304 nsew signal input
flabel metal2 s 601714 996690 601842 996890 0 FreeSans 320 90 0 0 gpio3_2_pad_a_esd_0_h
port 1305 nsew signal bidirectional
flabel metal2 s 600454 996690 600584 996890 0 FreeSans 320 90 0 0 gpio3_2_pad_a_esd_1_h
port 1306 nsew signal bidirectional
flabel metal2 s 599362 996690 599576 996890 0 FreeSans 320 90 0 0 gpio3_2_pad_a_noesd_h
port 1307 nsew signal bidirectional
flabel metal2 s 599058 996690 599110 996890 0 FreeSans 320 90 0 0 gpio3_2_analog_en
port 1308 nsew signal input
flabel metal2 s 596144 996690 596196 996890 0 FreeSans 320 90 0 0 gpio3_2_analog_pol
port 1309 nsew signal input
flabel metal2 s 595848 996690 595900 996890 0 FreeSans 320 90 0 0 gpio3_2_inp_dis
port 1310 nsew signal input
flabel metal2 s 594473 996690 594529 996890 0 FreeSans 320 90 0 0 gpio3_2_enable_inp_h
port 1311 nsew signal input
flabel metal2 s 593891 996690 593943 996890 0 FreeSans 320 90 0 0 gpio3_2_enable_h
port 1312 nsew signal input
flabel metal2 s 593162 996690 593214 996890 0 FreeSans 320 90 0 0 gpio3_2_hld_h_n
port 1313 nsew signal input
flabel metal2 s 592848 996690 592900 996890 0 FreeSans 320 90 0 0 gpio3_2_analog_sel
port 1314 nsew signal input
flabel metal2 s 592497 996690 592549 996890 0 FreeSans 320 90 0 0 gpio3_2_dm[2]
port 1315 nsew signal input
flabel metal2 s 600166 996690 600218 996890 0 FreeSans 320 90 0 0 gpio3_2_dm[1]
port 1316 nsew signal input
flabel metal2 s 596770 996690 596822 996890 0 FreeSans 320 90 0 0 gpio3_2_dm[0]
port 1317 nsew signal input
flabel metal2 s 592119 996690 592171 996890 0 FreeSans 320 90 0 0 gpio3_2_hld_ovr
port 1318 nsew signal input
flabel metal2 s 591270 996690 591322 996890 0 FreeSans 320 90 0 0 gpio3_2_out
port 1319 nsew signal input
flabel metal2 s 590061 996690 590113 996890 0 FreeSans 320 90 0 0 gpio3_2_enable_vswitch_h
port 1320 nsew signal input
flabel metal2 s 589350 996690 589402 996890 0 FreeSans 320 90 0 0 gpio3_2_enable_vdda_h
port 1321 nsew signal input
flabel metal2 s 588102 996690 588154 996890 0 FreeSans 320 90 0 0 gpio3_2_vtrip_sel
port 1322 nsew signal input
flabel metal2 s 587782 996690 587834 996890 0 FreeSans 320 90 0 0 gpio3_2_ib_mode_sel
port 1323 nsew signal input
flabel metal2 s 587468 996690 587520 996890 0 FreeSans 320 90 0 0 gpio3_2_oe_n
port 1324 nsew signal input
flabel metal2 s 586878 996690 587002 996890 0 FreeSans 320 90 0 0 gpio3_2_in_h
port 1325 nsew signal input
flabel metal2 s 604254 996690 604306 996890 0 FreeSans 320 90 0 0 gpio3_2_zero
port 1326 nsew signal output
flabel metal2 s 604616 996690 604668 996890 0 FreeSans 320 90 0 0 gpio3_2_one
port 1327 nsew signal output
flabel metal2 s 579290 996690 579342 996890 0 FreeSans 320 90 0 0 gpio3_3_tie_lo_esd
port 1328 nsew signal output
flabel metal2 s 578990 996690 579042 996890 0 FreeSans 320 90 0 0 gpio3_3_in
port 1329 nsew signal output
flabel metal2 s 578688 996690 578740 996890 0 FreeSans 320 90 0 0 gpio3_3_tie_hi_esd
port 1330 nsew signal output
flabel metal2 s 578390 996690 578442 996890 0 FreeSans 320 90 0 0 gpio3_3_enable_vddio
port 1331 nsew signal input
flabel metal2 s 578090 996690 578142 996890 0 FreeSans 320 90 0 0 gpio3_3_slow
port 1332 nsew signal input
flabel metal2 s 577714 996690 577842 996890 0 FreeSans 320 90 0 0 gpio3_3_pad_a_esd_0_h
port 1333 nsew signal bidirectional
flabel metal2 s 576454 996690 576584 996890 0 FreeSans 320 90 0 0 gpio3_3_pad_a_esd_1_h
port 1334 nsew signal bidirectional
flabel metal2 s 575362 996690 575576 996890 0 FreeSans 320 90 0 0 gpio3_3_pad_a_noesd_h
port 1335 nsew signal bidirectional
flabel metal2 s 575058 996690 575110 996890 0 FreeSans 320 90 0 0 gpio3_3_analog_en
port 1336 nsew signal input
flabel metal2 s 572144 996690 572196 996890 0 FreeSans 320 90 0 0 gpio3_3_analog_pol
port 1337 nsew signal input
flabel metal2 s 571848 996690 571900 996890 0 FreeSans 320 90 0 0 gpio3_3_inp_dis
port 1338 nsew signal input
flabel metal2 s 570473 996690 570529 996890 0 FreeSans 320 90 0 0 gpio3_3_enable_inp_h
port 1339 nsew signal input
flabel metal2 s 569891 996690 569943 996890 0 FreeSans 320 90 0 0 gpio3_3_enable_h
port 1340 nsew signal input
flabel metal2 s 569162 996690 569214 996890 0 FreeSans 320 90 0 0 gpio3_3_hld_h_n
port 1341 nsew signal input
flabel metal2 s 568848 996690 568900 996890 0 FreeSans 320 90 0 0 gpio3_3_analog_sel
port 1342 nsew signal input
flabel metal2 s 568497 996690 568549 996890 0 FreeSans 320 90 0 0 gpio3_3_dm[2]
port 1343 nsew signal input
flabel metal2 s 576166 996690 576218 996890 0 FreeSans 320 90 0 0 gpio3_3_dm[1]
port 1344 nsew signal input
flabel metal2 s 572770 996690 572822 996890 0 FreeSans 320 90 0 0 gpio3_3_dm[0]
port 1345 nsew signal input
flabel metal2 s 568119 996690 568171 996890 0 FreeSans 320 90 0 0 gpio3_3_hld_ovr
port 1346 nsew signal input
flabel metal2 s 567270 996690 567322 996890 0 FreeSans 320 90 0 0 gpio3_3_out
port 1347 nsew signal input
flabel metal2 s 566061 996690 566113 996890 0 FreeSans 320 90 0 0 gpio3_3_enable_vswitch_h
port 1348 nsew signal input
flabel metal2 s 565350 996690 565402 996890 0 FreeSans 320 90 0 0 gpio3_3_enable_vdda_h
port 1349 nsew signal input
flabel metal2 s 564102 996690 564154 996890 0 FreeSans 320 90 0 0 gpio3_3_vtrip_sel
port 1350 nsew signal input
flabel metal2 s 563782 996690 563834 996890 0 FreeSans 320 90 0 0 gpio3_3_ib_mode_sel
port 1351 nsew signal input
flabel metal2 s 563468 996690 563520 996890 0 FreeSans 320 90 0 0 gpio3_3_oe_n
port 1352 nsew signal input
flabel metal2 s 562878 996690 563002 996890 0 FreeSans 320 90 0 0 gpio3_3_in_h
port 1353 nsew signal input
flabel metal2 s 580254 996690 580306 996890 0 FreeSans 320 90 0 0 gpio3_3_zero
port 1354 nsew signal output
flabel metal2 s 580616 996690 580668 996890 0 FreeSans 320 90 0 0 gpio3_3_one
port 1355 nsew signal output
flabel metal2 s 509290 996690 509342 996890 0 FreeSans 320 90 0 0 gpio3_4_tie_lo_esd
port 1356 nsew signal output
flabel metal2 s 508990 996690 509042 996890 0 FreeSans 320 90 0 0 gpio3_4_in
port 1357 nsew signal output
flabel metal2 s 508688 996690 508740 996890 0 FreeSans 320 90 0 0 gpio3_4_tie_hi_esd
port 1358 nsew signal output
flabel metal2 s 508390 996690 508442 996890 0 FreeSans 320 90 0 0 gpio3_4_enable_vddio
port 1359 nsew signal input
flabel metal2 s 508090 996690 508142 996890 0 FreeSans 320 90 0 0 gpio3_4_slow
port 1360 nsew signal input
flabel metal2 s 507714 996690 507842 996890 0 FreeSans 320 90 0 0 gpio3_4_pad_a_esd_0_h
port 1361 nsew signal bidirectional
flabel metal2 s 506454 996690 506584 996890 0 FreeSans 320 90 0 0 gpio3_4_pad_a_esd_1_h
port 1362 nsew signal bidirectional
flabel metal2 s 505362 996690 505576 996890 0 FreeSans 320 90 0 0 gpio3_4_pad_a_noesd_h
port 1363 nsew signal bidirectional
flabel metal2 s 505058 996690 505110 996890 0 FreeSans 320 90 0 0 gpio3_4_analog_en
port 1364 nsew signal input
flabel metal2 s 502144 996690 502196 996890 0 FreeSans 320 90 0 0 gpio3_4_analog_pol
port 1365 nsew signal input
flabel metal2 s 501848 996690 501900 996890 0 FreeSans 320 90 0 0 gpio3_4_inp_dis
port 1366 nsew signal input
flabel metal2 s 500473 996690 500529 996890 0 FreeSans 320 90 0 0 gpio3_4_enable_inp_h
port 1367 nsew signal input
flabel metal2 s 499891 996690 499943 996890 0 FreeSans 320 90 0 0 gpio3_4_enable_h
port 1368 nsew signal input
flabel metal2 s 499162 996690 499214 996890 0 FreeSans 320 90 0 0 gpio3_4_hld_h_n
port 1369 nsew signal input
flabel metal2 s 498848 996690 498900 996890 0 FreeSans 320 90 0 0 gpio3_4_analog_sel
port 1370 nsew signal input
flabel metal2 s 498497 996690 498549 996890 0 FreeSans 320 90 0 0 gpio3_4_dm[2]
port 1371 nsew signal input
flabel metal2 s 506166 996690 506218 996890 0 FreeSans 320 90 0 0 gpio3_4_dm[1]
port 1372 nsew signal input
flabel metal2 s 502770 996690 502822 996890 0 FreeSans 320 90 0 0 gpio3_4_dm[0]
port 1373 nsew signal input
flabel metal2 s 498119 996690 498171 996890 0 FreeSans 320 90 0 0 gpio3_4_hld_ovr
port 1374 nsew signal input
flabel metal2 s 497270 996690 497322 996890 0 FreeSans 320 90 0 0 gpio3_4_out
port 1375 nsew signal input
flabel metal2 s 496061 996690 496113 996890 0 FreeSans 320 90 0 0 gpio3_4_enable_vswitch_h
port 1376 nsew signal input
flabel metal2 s 495350 996690 495402 996890 0 FreeSans 320 90 0 0 gpio3_4_enable_vdda_h
port 1377 nsew signal input
flabel metal2 s 494102 996690 494154 996890 0 FreeSans 320 90 0 0 gpio3_4_vtrip_sel
port 1378 nsew signal input
flabel metal2 s 493782 996690 493834 996890 0 FreeSans 320 90 0 0 gpio3_4_ib_mode_sel
port 1379 nsew signal input
flabel metal2 s 493468 996690 493520 996890 0 FreeSans 320 90 0 0 gpio3_4_oe_n
port 1380 nsew signal input
flabel metal2 s 492878 996690 493002 996890 0 FreeSans 320 90 0 0 gpio3_4_in_h
port 1381 nsew signal input
flabel metal2 s 510254 996690 510306 996890 0 FreeSans 320 90 0 0 gpio3_4_zero
port 1382 nsew signal output
flabel metal2 s 510616 996690 510668 996890 0 FreeSans 320 90 0 0 gpio3_4_one
port 1383 nsew signal output
flabel metal2 s 485290 996690 485342 996890 0 FreeSans 320 90 0 0 gpio3_5_tie_lo_esd
port 1384 nsew signal output
flabel metal2 s 484990 996690 485042 996890 0 FreeSans 320 90 0 0 gpio3_5_in
port 1385 nsew signal output
flabel metal2 s 484688 996690 484740 996890 0 FreeSans 320 90 0 0 gpio3_5_tie_hi_esd
port 1386 nsew signal output
flabel metal2 s 484390 996690 484442 996890 0 FreeSans 320 90 0 0 gpio3_5_enable_vddio
port 1387 nsew signal input
flabel metal2 s 484090 996690 484142 996890 0 FreeSans 320 90 0 0 gpio3_5_slow
port 1388 nsew signal input
flabel metal2 s 483714 996690 483842 996890 0 FreeSans 320 90 0 0 gpio3_5_pad_a_esd_0_h
port 1389 nsew signal bidirectional
flabel metal2 s 482454 996690 482584 996890 0 FreeSans 320 90 0 0 gpio3_5_pad_a_esd_1_h
port 1390 nsew signal bidirectional
flabel metal2 s 481362 996690 481576 996890 0 FreeSans 320 90 0 0 gpio3_5_pad_a_noesd_h
port 1391 nsew signal bidirectional
flabel metal2 s 481058 996690 481110 996890 0 FreeSans 320 90 0 0 gpio3_5_analog_en
port 1392 nsew signal input
flabel metal2 s 478144 996690 478196 996890 0 FreeSans 320 90 0 0 gpio3_5_analog_pol
port 1393 nsew signal input
flabel metal2 s 477848 996690 477900 996890 0 FreeSans 320 90 0 0 gpio3_5_inp_dis
port 1394 nsew signal input
flabel metal2 s 476473 996690 476529 996890 0 FreeSans 320 90 0 0 gpio3_5_enable_inp_h
port 1395 nsew signal input
flabel metal2 s 475891 996690 475943 996890 0 FreeSans 320 90 0 0 gpio3_5_enable_h
port 1396 nsew signal input
flabel metal2 s 475162 996690 475214 996890 0 FreeSans 320 90 0 0 gpio3_5_hld_h_n
port 1397 nsew signal input
flabel metal2 s 474848 996690 474900 996890 0 FreeSans 320 90 0 0 gpio3_5_analog_sel
port 1398 nsew signal input
flabel metal2 s 474497 996690 474549 996890 0 FreeSans 320 90 0 0 gpio3_5_dm[2]
port 1399 nsew signal input
flabel metal2 s 482166 996690 482218 996890 0 FreeSans 320 90 0 0 gpio3_5_dm[1]
port 1400 nsew signal input
flabel metal2 s 478770 996690 478822 996890 0 FreeSans 320 90 0 0 gpio3_5_dm[0]
port 1401 nsew signal input
flabel metal2 s 474119 996690 474171 996890 0 FreeSans 320 90 0 0 gpio3_5_hld_ovr
port 1402 nsew signal input
flabel metal2 s 473270 996690 473322 996890 0 FreeSans 320 90 0 0 gpio3_5_out
port 1403 nsew signal input
flabel metal2 s 472061 996690 472113 996890 0 FreeSans 320 90 0 0 gpio3_5_enable_vswitch_h
port 1404 nsew signal input
flabel metal2 s 471350 996690 471402 996890 0 FreeSans 320 90 0 0 gpio3_5_enable_vdda_h
port 1405 nsew signal input
flabel metal2 s 470102 996690 470154 996890 0 FreeSans 320 90 0 0 gpio3_5_vtrip_sel
port 1406 nsew signal input
flabel metal2 s 469782 996690 469834 996890 0 FreeSans 320 90 0 0 gpio3_5_ib_mode_sel
port 1407 nsew signal input
flabel metal2 s 469468 996690 469520 996890 0 FreeSans 320 90 0 0 gpio3_5_oe_n
port 1408 nsew signal input
flabel metal2 s 468878 996690 469002 996890 0 FreeSans 320 90 0 0 gpio3_5_in_h
port 1409 nsew signal input
flabel metal2 s 486254 996690 486306 996890 0 FreeSans 320 90 0 0 gpio3_5_zero
port 1410 nsew signal output
flabel metal2 s 486616 996690 486668 996890 0 FreeSans 320 90 0 0 gpio3_5_one
port 1411 nsew signal output
flabel metal2 s 461290 996690 461342 996890 0 FreeSans 320 90 0 0 gpio3_6_tie_lo_esd
port 1412 nsew signal output
flabel metal2 s 460990 996690 461042 996890 0 FreeSans 320 90 0 0 gpio3_6_in
port 1413 nsew signal output
flabel metal2 s 460688 996690 460740 996890 0 FreeSans 320 90 0 0 gpio3_6_tie_hi_esd
port 1414 nsew signal output
flabel metal2 s 460390 996690 460442 996890 0 FreeSans 320 90 0 0 gpio3_6_enable_vddio
port 1415 nsew signal input
flabel metal2 s 460090 996690 460142 996890 0 FreeSans 320 90 0 0 gpio3_6_slow
port 1416 nsew signal input
flabel metal2 s 459714 996690 459842 996890 0 FreeSans 320 90 0 0 gpio3_6_pad_a_esd_0_h
port 1417 nsew signal bidirectional
flabel metal2 s 458454 996690 458584 996890 0 FreeSans 320 90 0 0 gpio3_6_pad_a_esd_1_h
port 1418 nsew signal bidirectional
flabel metal2 s 457362 996690 457576 996890 0 FreeSans 320 90 0 0 gpio3_6_pad_a_noesd_h
port 1419 nsew signal bidirectional
flabel metal2 s 457058 996690 457110 996890 0 FreeSans 320 90 0 0 gpio3_6_analog_en
port 1420 nsew signal input
flabel metal2 s 454144 996690 454196 996890 0 FreeSans 320 90 0 0 gpio3_6_analog_pol
port 1421 nsew signal input
flabel metal2 s 453848 996690 453900 996890 0 FreeSans 320 90 0 0 gpio3_6_inp_dis
port 1422 nsew signal input
flabel metal2 s 452473 996690 452529 996890 0 FreeSans 320 90 0 0 gpio3_6_enable_inp_h
port 1423 nsew signal input
flabel metal2 s 451891 996690 451943 996890 0 FreeSans 320 90 0 0 gpio3_6_enable_h
port 1424 nsew signal input
flabel metal2 s 451162 996690 451214 996890 0 FreeSans 320 90 0 0 gpio3_6_hld_h_n
port 1425 nsew signal input
flabel metal2 s 450848 996690 450900 996890 0 FreeSans 320 90 0 0 gpio3_6_analog_sel
port 1426 nsew signal input
flabel metal2 s 450497 996690 450549 996890 0 FreeSans 320 90 0 0 gpio3_6_dm[2]
port 1427 nsew signal input
flabel metal2 s 458166 996690 458218 996890 0 FreeSans 320 90 0 0 gpio3_6_dm[1]
port 1428 nsew signal input
flabel metal2 s 454770 996690 454822 996890 0 FreeSans 320 90 0 0 gpio3_6_dm[0]
port 1429 nsew signal input
flabel metal2 s 450119 996690 450171 996890 0 FreeSans 320 90 0 0 gpio3_6_hld_ovr
port 1430 nsew signal input
flabel metal2 s 449270 996690 449322 996890 0 FreeSans 320 90 0 0 gpio3_6_out
port 1431 nsew signal input
flabel metal2 s 448061 996690 448113 996890 0 FreeSans 320 90 0 0 gpio3_6_enable_vswitch_h
port 1432 nsew signal input
flabel metal2 s 447350 996690 447402 996890 0 FreeSans 320 90 0 0 gpio3_6_enable_vdda_h
port 1433 nsew signal input
flabel metal2 s 446102 996690 446154 996890 0 FreeSans 320 90 0 0 gpio3_6_vtrip_sel
port 1434 nsew signal input
flabel metal2 s 445782 996690 445834 996890 0 FreeSans 320 90 0 0 gpio3_6_ib_mode_sel
port 1435 nsew signal input
flabel metal2 s 445468 996690 445520 996890 0 FreeSans 320 90 0 0 gpio3_6_oe_n
port 1436 nsew signal input
flabel metal2 s 444878 996690 445002 996890 0 FreeSans 320 90 0 0 gpio3_6_in_h
port 1437 nsew signal input
flabel metal2 s 462254 996690 462306 996890 0 FreeSans 320 90 0 0 gpio3_6_zero
port 1438 nsew signal output
flabel metal2 s 462616 996690 462668 996890 0 FreeSans 320 90 0 0 gpio3_6_one
port 1439 nsew signal output
flabel metal2 s 437290 996690 437342 996890 0 FreeSans 320 90 0 0 gpio3_7_tie_lo_esd
port 1440 nsew signal output
flabel metal2 s 436990 996690 437042 996890 0 FreeSans 320 90 0 0 gpio3_7_in
port 1441 nsew signal output
flabel metal2 s 436688 996690 436740 996890 0 FreeSans 320 90 0 0 gpio3_7_tie_hi_esd
port 1442 nsew signal output
flabel metal2 s 436390 996690 436442 996890 0 FreeSans 320 90 0 0 gpio3_7_enable_vddio
port 1443 nsew signal input
flabel metal2 s 436090 996690 436142 996890 0 FreeSans 320 90 0 0 gpio3_7_slow
port 1444 nsew signal input
flabel metal2 s 435714 996690 435842 996890 0 FreeSans 320 90 0 0 gpio3_7_pad_a_esd_0_h
port 1445 nsew signal bidirectional
flabel metal2 s 434454 996690 434584 996890 0 FreeSans 320 90 0 0 gpio3_7_pad_a_esd_1_h
port 1446 nsew signal bidirectional
flabel metal2 s 433362 996690 433576 996890 0 FreeSans 320 90 0 0 gpio3_7_pad_a_noesd_h
port 1447 nsew signal bidirectional
flabel metal2 s 433058 996690 433110 996890 0 FreeSans 320 90 0 0 gpio3_7_analog_en
port 1448 nsew signal input
flabel metal2 s 430144 996690 430196 996890 0 FreeSans 320 90 0 0 gpio3_7_analog_pol
port 1449 nsew signal input
flabel metal2 s 429848 996690 429900 996890 0 FreeSans 320 90 0 0 gpio3_7_inp_dis
port 1450 nsew signal input
flabel metal2 s 428473 996690 428529 996890 0 FreeSans 320 90 0 0 gpio3_7_enable_inp_h
port 1451 nsew signal input
flabel metal2 s 427891 996690 427943 996890 0 FreeSans 320 90 0 0 gpio3_7_enable_h
port 1452 nsew signal input
flabel metal2 s 427162 996690 427214 996890 0 FreeSans 320 90 0 0 gpio3_7_hld_h_n
port 1453 nsew signal input
flabel metal2 s 426848 996690 426900 996890 0 FreeSans 320 90 0 0 gpio3_7_analog_sel
port 1454 nsew signal input
flabel metal2 s 426497 996690 426549 996890 0 FreeSans 320 90 0 0 gpio3_7_dm[2]
port 1455 nsew signal input
flabel metal2 s 434166 996690 434218 996890 0 FreeSans 320 90 0 0 gpio3_7_dm[1]
port 1456 nsew signal input
flabel metal2 s 430770 996690 430822 996890 0 FreeSans 320 90 0 0 gpio3_7_dm[0]
port 1457 nsew signal input
flabel metal2 s 426119 996690 426171 996890 0 FreeSans 320 90 0 0 gpio3_7_hld_ovr
port 1458 nsew signal input
flabel metal2 s 425270 996690 425322 996890 0 FreeSans 320 90 0 0 gpio3_7_out
port 1459 nsew signal input
flabel metal2 s 424061 996690 424113 996890 0 FreeSans 320 90 0 0 gpio3_7_enable_vswitch_h
port 1460 nsew signal input
flabel metal2 s 423350 996690 423402 996890 0 FreeSans 320 90 0 0 gpio3_7_enable_vdda_h
port 1461 nsew signal input
flabel metal2 s 422102 996690 422154 996890 0 FreeSans 320 90 0 0 gpio3_7_vtrip_sel
port 1462 nsew signal input
flabel metal2 s 421782 996690 421834 996890 0 FreeSans 320 90 0 0 gpio3_7_ib_mode_sel
port 1463 nsew signal input
flabel metal2 s 421468 996690 421520 996890 0 FreeSans 320 90 0 0 gpio3_7_oe_n
port 1464 nsew signal input
flabel metal2 s 420878 996690 421002 996890 0 FreeSans 320 90 0 0 gpio3_7_in_h
port 1465 nsew signal input
flabel metal2 s 438254 996690 438306 996890 0 FreeSans 320 90 0 0 gpio3_7_zero
port 1466 nsew signal output
flabel metal2 s 438616 996690 438668 996890 0 FreeSans 320 90 0 0 gpio3_7_one
port 1467 nsew signal output
flabel metal2 s 359566 996600 361362 997000 0 FreeSans 320 0 0 0 analog_0_core
port 1468 nsew analog bidirectional
flabel metal2 s 336566 996600 338362 997000 0 FreeSans 320 0 0 0 analog_1_core
port 1469 nsew analog bidirectional
flabel metal2 s 298290 996690 298342 996890 0 FreeSans 320 90 0 0 gpio4_0_tie_lo_esd
port 1470 nsew signal output
flabel metal2 s 297990 996690 298042 996890 0 FreeSans 320 90 0 0 gpio4_0_in
port 1471 nsew signal output
flabel metal2 s 297688 996690 297740 996890 0 FreeSans 320 90 0 0 gpio4_0_tie_hi_esd
port 1472 nsew signal output
flabel metal2 s 297390 996690 297442 996890 0 FreeSans 320 90 0 0 gpio4_0_enable_vddio
port 1473 nsew signal input
flabel metal2 s 297090 996690 297142 996890 0 FreeSans 320 90 0 0 gpio4_0_slow
port 1474 nsew signal input
flabel metal2 s 296714 996690 296842 996890 0 FreeSans 320 90 0 0 gpio4_0_pad_a_esd_0_h
port 1475 nsew signal bidirectional
flabel metal2 s 295454 996690 295584 996890 0 FreeSans 320 90 0 0 gpio4_0_pad_a_esd_1_h
port 1476 nsew signal bidirectional
flabel metal2 s 294362 996690 294576 996890 0 FreeSans 320 90 0 0 gpio4_0_pad_a_noesd_h
port 1477 nsew signal bidirectional
flabel metal2 s 294058 996690 294110 996890 0 FreeSans 320 90 0 0 gpio4_0_analog_en
port 1478 nsew signal input
flabel metal2 s 291144 996690 291196 996890 0 FreeSans 320 90 0 0 gpio4_0_analog_pol
port 1479 nsew signal input
flabel metal2 s 290848 996690 290900 996890 0 FreeSans 320 90 0 0 gpio4_0_inp_dis
port 1480 nsew signal input
flabel metal2 s 289473 996690 289529 996890 0 FreeSans 320 90 0 0 gpio4_0_enable_inp_h
port 1481 nsew signal input
flabel metal2 s 288891 996690 288943 996890 0 FreeSans 320 90 0 0 gpio4_0_enable_h
port 1482 nsew signal input
flabel metal2 s 288162 996690 288214 996890 0 FreeSans 320 90 0 0 gpio4_0_hld_h_n
port 1483 nsew signal input
flabel metal2 s 287848 996690 287900 996890 0 FreeSans 320 90 0 0 gpio4_0_analog_sel
port 1484 nsew signal input
flabel metal2 s 287497 996690 287549 996890 0 FreeSans 320 90 0 0 gpio4_0_dm[2]
port 1485 nsew signal input
flabel metal2 s 295166 996690 295218 996890 0 FreeSans 320 90 0 0 gpio4_0_dm[1]
port 1486 nsew signal input
flabel metal2 s 291770 996690 291822 996890 0 FreeSans 320 90 0 0 gpio4_0_dm[0]
port 1487 nsew signal input
flabel metal2 s 287119 996690 287171 996890 0 FreeSans 320 90 0 0 gpio4_0_hld_ovr
port 1488 nsew signal input
flabel metal2 s 286270 996690 286322 996890 0 FreeSans 320 90 0 0 gpio4_0_out
port 1489 nsew signal input
flabel metal2 s 285061 996690 285113 996890 0 FreeSans 320 90 0 0 gpio4_0_enable_vswitch_h
port 1490 nsew signal input
flabel metal2 s 284350 996690 284402 996890 0 FreeSans 320 90 0 0 gpio4_0_enable_vdda_h
port 1491 nsew signal input
flabel metal2 s 283102 996690 283154 996890 0 FreeSans 320 90 0 0 gpio4_0_vtrip_sel
port 1492 nsew signal input
flabel metal2 s 282782 996690 282834 996890 0 FreeSans 320 90 0 0 gpio4_0_ib_mode_sel
port 1493 nsew signal input
flabel metal2 s 282468 996690 282520 996890 0 FreeSans 320 90 0 0 gpio4_0_oe_n
port 1494 nsew signal input
flabel metal2 s 281878 996690 282002 996890 0 FreeSans 320 90 0 0 gpio4_0_in_h
port 1495 nsew signal input
flabel metal2 s 299254 996690 299306 996890 0 FreeSans 320 90 0 0 gpio4_0_zero
port 1496 nsew signal output
flabel metal2 s 299616 996690 299668 996890 0 FreeSans 320 90 0 0 gpio4_0_one
port 1497 nsew signal output
flabel metal2 s 274290 996690 274342 996890 0 FreeSans 320 90 0 0 gpio4_1_tie_lo_esd
port 1498 nsew signal output
flabel metal2 s 273990 996690 274042 996890 0 FreeSans 320 90 0 0 gpio4_1_in
port 1499 nsew signal output
flabel metal2 s 273688 996690 273740 996890 0 FreeSans 320 90 0 0 gpio4_1_tie_hi_esd
port 1500 nsew signal output
flabel metal2 s 273390 996690 273442 996890 0 FreeSans 320 90 0 0 gpio4_1_enable_vddio
port 1501 nsew signal input
flabel metal2 s 273090 996690 273142 996890 0 FreeSans 320 90 0 0 gpio4_1_slow
port 1502 nsew signal input
flabel metal2 s 272714 996690 272842 996890 0 FreeSans 320 90 0 0 gpio4_1_pad_a_esd_0_h
port 1503 nsew signal bidirectional
flabel metal2 s 271454 996690 271584 996890 0 FreeSans 320 90 0 0 gpio4_1_pad_a_esd_1_h
port 1504 nsew signal bidirectional
flabel metal2 s 270362 996690 270576 996890 0 FreeSans 320 90 0 0 gpio4_1_pad_a_noesd_h
port 1505 nsew signal bidirectional
flabel metal2 s 270058 996690 270110 996890 0 FreeSans 320 90 0 0 gpio4_1_analog_en
port 1506 nsew signal input
flabel metal2 s 267144 996690 267196 996890 0 FreeSans 320 90 0 0 gpio4_1_analog_pol
port 1507 nsew signal input
flabel metal2 s 266848 996690 266900 996890 0 FreeSans 320 90 0 0 gpio4_1_inp_dis
port 1508 nsew signal input
flabel metal2 s 265473 996690 265529 996890 0 FreeSans 320 90 0 0 gpio4_1_enable_inp_h
port 1509 nsew signal input
flabel metal2 s 264891 996690 264943 996890 0 FreeSans 320 90 0 0 gpio4_1_enable_h
port 1510 nsew signal input
flabel metal2 s 264162 996690 264214 996890 0 FreeSans 320 90 0 0 gpio4_1_hld_h_n
port 1511 nsew signal input
flabel metal2 s 263848 996690 263900 996890 0 FreeSans 320 90 0 0 gpio4_1_analog_sel
port 1512 nsew signal input
flabel metal2 s 263497 996690 263549 996890 0 FreeSans 320 90 0 0 gpio4_1_dm[2]
port 1513 nsew signal input
flabel metal2 s 271166 996690 271218 996890 0 FreeSans 320 90 0 0 gpio4_1_dm[1]
port 1514 nsew signal input
flabel metal2 s 267770 996690 267822 996890 0 FreeSans 320 90 0 0 gpio4_1_dm[0]
port 1515 nsew signal input
flabel metal2 s 263119 996690 263171 996890 0 FreeSans 320 90 0 0 gpio4_1_hld_ovr
port 1516 nsew signal input
flabel metal2 s 262270 996690 262322 996890 0 FreeSans 320 90 0 0 gpio4_1_out
port 1517 nsew signal input
flabel metal2 s 261061 996690 261113 996890 0 FreeSans 320 90 0 0 gpio4_1_enable_vswitch_h
port 1518 nsew signal input
flabel metal2 s 260350 996690 260402 996890 0 FreeSans 320 90 0 0 gpio4_1_enable_vdda_h
port 1519 nsew signal input
flabel metal2 s 259102 996690 259154 996890 0 FreeSans 320 90 0 0 gpio4_1_vtrip_sel
port 1520 nsew signal input
flabel metal2 s 258782 996690 258834 996890 0 FreeSans 320 90 0 0 gpio4_1_ib_mode_sel
port 1521 nsew signal input
flabel metal2 s 258468 996690 258520 996890 0 FreeSans 320 90 0 0 gpio4_1_oe_n
port 1522 nsew signal input
flabel metal2 s 257878 996690 258002 996890 0 FreeSans 320 90 0 0 gpio4_1_in_h
port 1523 nsew signal input
flabel metal2 s 275254 996690 275306 996890 0 FreeSans 320 90 0 0 gpio4_1_zero
port 1524 nsew signal output
flabel metal2 s 275616 996690 275668 996890 0 FreeSans 320 90 0 0 gpio4_1_one
port 1525 nsew signal output
flabel metal2 s 250290 996690 250342 996890 0 FreeSans 320 90 0 0 gpio4_2_tie_lo_esd
port 1526 nsew signal output
flabel metal2 s 249990 996690 250042 996890 0 FreeSans 320 90 0 0 gpio4_2_in
port 1527 nsew signal output
flabel metal2 s 249688 996690 249740 996890 0 FreeSans 320 90 0 0 gpio4_2_tie_hi_esd
port 1528 nsew signal output
flabel metal2 s 249390 996690 249442 996890 0 FreeSans 320 90 0 0 gpio4_2_enable_vddio
port 1529 nsew signal input
flabel metal2 s 249090 996690 249142 996890 0 FreeSans 320 90 0 0 gpio4_2_slow
port 1530 nsew signal input
flabel metal2 s 248714 996690 248842 996890 0 FreeSans 320 90 0 0 gpio4_2_pad_a_esd_0_h
port 1531 nsew signal bidirectional
flabel metal2 s 247454 996690 247584 996890 0 FreeSans 320 90 0 0 gpio4_2_pad_a_esd_1_h
port 1532 nsew signal bidirectional
flabel metal2 s 246362 996690 246576 996890 0 FreeSans 320 90 0 0 gpio4_2_pad_a_noesd_h
port 1533 nsew signal bidirectional
flabel metal2 s 246058 996690 246110 996890 0 FreeSans 320 90 0 0 gpio4_2_analog_en
port 1534 nsew signal input
flabel metal2 s 243144 996690 243196 996890 0 FreeSans 320 90 0 0 gpio4_2_analog_pol
port 1535 nsew signal input
flabel metal2 s 242848 996690 242900 996890 0 FreeSans 320 90 0 0 gpio4_2_inp_dis
port 1536 nsew signal input
flabel metal2 s 241473 996690 241529 996890 0 FreeSans 320 90 0 0 gpio4_2_enable_inp_h
port 1537 nsew signal input
flabel metal2 s 240891 996690 240943 996890 0 FreeSans 320 90 0 0 gpio4_2_enable_h
port 1538 nsew signal input
flabel metal2 s 240162 996690 240214 996890 0 FreeSans 320 90 0 0 gpio4_2_hld_h_n
port 1539 nsew signal input
flabel metal2 s 239848 996690 239900 996890 0 FreeSans 320 90 0 0 gpio4_2_analog_sel
port 1540 nsew signal input
flabel metal2 s 239497 996690 239549 996890 0 FreeSans 320 90 0 0 gpio4_2_dm[2]
port 1541 nsew signal input
flabel metal2 s 247166 996690 247218 996890 0 FreeSans 320 90 0 0 gpio4_2_dm[1]
port 1542 nsew signal input
flabel metal2 s 243770 996690 243822 996890 0 FreeSans 320 90 0 0 gpio4_2_dm[0]
port 1543 nsew signal input
flabel metal2 s 239119 996690 239171 996890 0 FreeSans 320 90 0 0 gpio4_2_hld_ovr
port 1544 nsew signal input
flabel metal2 s 238270 996690 238322 996890 0 FreeSans 320 90 0 0 gpio4_2_out
port 1545 nsew signal input
flabel metal2 s 237061 996690 237113 996890 0 FreeSans 320 90 0 0 gpio4_2_enable_vswitch_h
port 1546 nsew signal input
flabel metal2 s 236350 996690 236402 996890 0 FreeSans 320 90 0 0 gpio4_2_enable_vdda_h
port 1547 nsew signal input
flabel metal2 s 235102 996690 235154 996890 0 FreeSans 320 90 0 0 gpio4_2_vtrip_sel
port 1548 nsew signal input
flabel metal2 s 234782 996690 234834 996890 0 FreeSans 320 90 0 0 gpio4_2_ib_mode_sel
port 1549 nsew signal input
flabel metal2 s 234468 996690 234520 996890 0 FreeSans 320 90 0 0 gpio4_2_oe_n
port 1550 nsew signal input
flabel metal2 s 233878 996690 234002 996890 0 FreeSans 320 90 0 0 gpio4_2_in_h
port 1551 nsew signal input
flabel metal2 s 251254 996690 251306 996890 0 FreeSans 320 90 0 0 gpio4_2_zero
port 1552 nsew signal output
flabel metal2 s 251616 996690 251668 996890 0 FreeSans 320 90 0 0 gpio4_2_one
port 1553 nsew signal output
flabel metal2 s 226290 996690 226342 996890 0 FreeSans 320 90 0 0 gpio4_3_tie_lo_esd
port 1554 nsew signal output
flabel metal2 s 225990 996690 226042 996890 0 FreeSans 320 90 0 0 gpio4_3_in
port 1555 nsew signal output
flabel metal2 s 225688 996690 225740 996890 0 FreeSans 320 90 0 0 gpio4_3_tie_hi_esd
port 1556 nsew signal output
flabel metal2 s 225390 996690 225442 996890 0 FreeSans 320 90 0 0 gpio4_3_enable_vddio
port 1557 nsew signal input
flabel metal2 s 225090 996690 225142 996890 0 FreeSans 320 90 0 0 gpio4_3_slow
port 1558 nsew signal input
flabel metal2 s 224714 996690 224842 996890 0 FreeSans 320 90 0 0 gpio4_3_pad_a_esd_0_h
port 1559 nsew signal bidirectional
flabel metal2 s 223454 996690 223584 996890 0 FreeSans 320 90 0 0 gpio4_3_pad_a_esd_1_h
port 1560 nsew signal bidirectional
flabel metal2 s 222362 996690 222576 996890 0 FreeSans 320 90 0 0 gpio4_3_pad_a_noesd_h
port 1561 nsew signal bidirectional
flabel metal2 s 222058 996690 222110 996890 0 FreeSans 320 90 0 0 gpio4_3_analog_en
port 1562 nsew signal input
flabel metal2 s 219144 996690 219196 996890 0 FreeSans 320 90 0 0 gpio4_3_analog_pol
port 1563 nsew signal input
flabel metal2 s 218848 996690 218900 996890 0 FreeSans 320 90 0 0 gpio4_3_inp_dis
port 1564 nsew signal input
flabel metal2 s 217473 996690 217529 996890 0 FreeSans 320 90 0 0 gpio4_3_enable_inp_h
port 1565 nsew signal input
flabel metal2 s 216891 996690 216943 996890 0 FreeSans 320 90 0 0 gpio4_3_enable_h
port 1566 nsew signal input
flabel metal2 s 216162 996690 216214 996890 0 FreeSans 320 90 0 0 gpio4_3_hld_h_n
port 1567 nsew signal input
flabel metal2 s 215848 996690 215900 996890 0 FreeSans 320 90 0 0 gpio4_3_analog_sel
port 1568 nsew signal input
flabel metal2 s 215497 996690 215549 996890 0 FreeSans 320 90 0 0 gpio4_3_dm[2]
port 1569 nsew signal input
flabel metal2 s 223166 996690 223218 996890 0 FreeSans 320 90 0 0 gpio4_3_dm[1]
port 1570 nsew signal input
flabel metal2 s 219770 996690 219822 996890 0 FreeSans 320 90 0 0 gpio4_3_dm[0]
port 1571 nsew signal input
flabel metal2 s 215119 996690 215171 996890 0 FreeSans 320 90 0 0 gpio4_3_hld_ovr
port 1572 nsew signal input
flabel metal2 s 214270 996690 214322 996890 0 FreeSans 320 90 0 0 gpio4_3_out
port 1573 nsew signal input
flabel metal2 s 213061 996690 213113 996890 0 FreeSans 320 90 0 0 gpio4_3_enable_vswitch_h
port 1574 nsew signal input
flabel metal2 s 212350 996690 212402 996890 0 FreeSans 320 90 0 0 gpio4_3_enable_vdda_h
port 1575 nsew signal input
flabel metal2 s 211102 996690 211154 996890 0 FreeSans 320 90 0 0 gpio4_3_vtrip_sel
port 1576 nsew signal input
flabel metal2 s 210782 996690 210834 996890 0 FreeSans 320 90 0 0 gpio4_3_ib_mode_sel
port 1577 nsew signal input
flabel metal2 s 210468 996690 210520 996890 0 FreeSans 320 90 0 0 gpio4_3_oe_n
port 1578 nsew signal input
flabel metal2 s 209878 996690 210002 996890 0 FreeSans 320 90 0 0 gpio4_3_in_h
port 1579 nsew signal input
flabel metal2 s 227254 996690 227306 996890 0 FreeSans 320 90 0 0 gpio4_3_zero
port 1580 nsew signal output
flabel metal2 s 227616 996690 227668 996890 0 FreeSans 320 90 0 0 gpio4_3_one
port 1581 nsew signal output
flabel metal2 s 156290 996690 156342 996890 0 FreeSans 320 90 0 0 gpio4_4_tie_lo_esd
port 1582 nsew signal output
flabel metal2 s 155990 996690 156042 996890 0 FreeSans 320 90 0 0 gpio4_4_in
port 1583 nsew signal output
flabel metal2 s 155688 996690 155740 996890 0 FreeSans 320 90 0 0 gpio4_4_tie_hi_esd
port 1584 nsew signal output
flabel metal2 s 155390 996690 155442 996890 0 FreeSans 320 90 0 0 gpio4_4_enable_vddio
port 1585 nsew signal input
flabel metal2 s 155090 996690 155142 996890 0 FreeSans 320 90 0 0 gpio4_4_slow
port 1586 nsew signal input
flabel metal2 s 154714 996690 154842 996890 0 FreeSans 320 90 0 0 gpio4_4_pad_a_esd_0_h
port 1587 nsew signal bidirectional
flabel metal2 s 153454 996690 153584 996890 0 FreeSans 320 90 0 0 gpio4_4_pad_a_esd_1_h
port 1588 nsew signal bidirectional
flabel metal2 s 152362 996690 152576 996890 0 FreeSans 320 90 0 0 gpio4_4_pad_a_noesd_h
port 1589 nsew signal bidirectional
flabel metal2 s 152058 996690 152110 996890 0 FreeSans 320 90 0 0 gpio4_4_analog_en
port 1590 nsew signal input
flabel metal2 s 149144 996690 149196 996890 0 FreeSans 320 90 0 0 gpio4_4_analog_pol
port 1591 nsew signal input
flabel metal2 s 148848 996690 148900 996890 0 FreeSans 320 90 0 0 gpio4_4_inp_dis
port 1592 nsew signal input
flabel metal2 s 147473 996690 147529 996890 0 FreeSans 320 90 0 0 gpio4_4_enable_inp_h
port 1593 nsew signal input
flabel metal2 s 146891 996690 146943 996890 0 FreeSans 320 90 0 0 gpio4_4_enable_h
port 1594 nsew signal input
flabel metal2 s 146162 996690 146214 996890 0 FreeSans 320 90 0 0 gpio4_4_hld_h_n
port 1595 nsew signal input
flabel metal2 s 145848 996690 145900 996890 0 FreeSans 320 90 0 0 gpio4_4_analog_sel
port 1596 nsew signal input
flabel metal2 s 145497 996690 145549 996890 0 FreeSans 320 90 0 0 gpio4_4_dm[2]
port 1597 nsew signal input
flabel metal2 s 153166 996690 153218 996890 0 FreeSans 320 90 0 0 gpio4_4_dm[1]
port 1598 nsew signal input
flabel metal2 s 149770 996690 149822 996890 0 FreeSans 320 90 0 0 gpio4_4_dm[0]
port 1599 nsew signal input
flabel metal2 s 145119 996690 145171 996890 0 FreeSans 320 90 0 0 gpio4_4_hld_ovr
port 1600 nsew signal input
flabel metal2 s 144270 996690 144322 996890 0 FreeSans 320 90 0 0 gpio4_4_out
port 1601 nsew signal input
flabel metal2 s 143061 996690 143113 996890 0 FreeSans 320 90 0 0 gpio4_4_enable_vswitch_h
port 1602 nsew signal input
flabel metal2 s 142350 996690 142402 996890 0 FreeSans 320 90 0 0 gpio4_4_enable_vdda_h
port 1603 nsew signal input
flabel metal2 s 141102 996690 141154 996890 0 FreeSans 320 90 0 0 gpio4_4_vtrip_sel
port 1604 nsew signal input
flabel metal2 s 140782 996690 140834 996890 0 FreeSans 320 90 0 0 gpio4_4_ib_mode_sel
port 1605 nsew signal input
flabel metal2 s 140468 996690 140520 996890 0 FreeSans 320 90 0 0 gpio4_4_oe_n
port 1606 nsew signal input
flabel metal2 s 139878 996690 140002 996890 0 FreeSans 320 90 0 0 gpio4_4_in_h
port 1607 nsew signal input
flabel metal2 s 157254 996690 157306 996890 0 FreeSans 320 90 0 0 gpio4_4_zero
port 1608 nsew signal output
flabel metal2 s 157616 996690 157668 996890 0 FreeSans 320 90 0 0 gpio4_4_one
port 1609 nsew signal output
flabel metal2 s 132290 996690 132342 996890 0 FreeSans 320 90 0 0 gpio4_5_tie_lo_esd
port 1610 nsew signal output
flabel metal2 s 131990 996690 132042 996890 0 FreeSans 320 90 0 0 gpio4_5_in
port 1611 nsew signal output
flabel metal2 s 131688 996690 131740 996890 0 FreeSans 320 90 0 0 gpio4_5_tie_hi_esd
port 1612 nsew signal output
flabel metal2 s 131390 996690 131442 996890 0 FreeSans 320 90 0 0 gpio4_5_enable_vddio
port 1613 nsew signal input
flabel metal2 s 131090 996690 131142 996890 0 FreeSans 320 90 0 0 gpio4_5_slow
port 1614 nsew signal input
flabel metal2 s 130714 996690 130842 996890 0 FreeSans 320 90 0 0 gpio4_5_pad_a_esd_0_h
port 1615 nsew signal bidirectional
flabel metal2 s 129454 996690 129584 996890 0 FreeSans 320 90 0 0 gpio4_5_pad_a_esd_1_h
port 1616 nsew signal bidirectional
flabel metal2 s 128362 996690 128576 996890 0 FreeSans 320 90 0 0 gpio4_5_pad_a_noesd_h
port 1617 nsew signal bidirectional
flabel metal2 s 128058 996690 128110 996890 0 FreeSans 320 90 0 0 gpio4_5_analog_en
port 1618 nsew signal input
flabel metal2 s 125144 996690 125196 996890 0 FreeSans 320 90 0 0 gpio4_5_analog_pol
port 1619 nsew signal input
flabel metal2 s 124848 996690 124900 996890 0 FreeSans 320 90 0 0 gpio4_5_inp_dis
port 1620 nsew signal input
flabel metal2 s 123473 996690 123529 996890 0 FreeSans 320 90 0 0 gpio4_5_enable_inp_h
port 1621 nsew signal input
flabel metal2 s 122891 996690 122943 996890 0 FreeSans 320 90 0 0 gpio4_5_enable_h
port 1622 nsew signal input
flabel metal2 s 122162 996690 122214 996890 0 FreeSans 320 90 0 0 gpio4_5_hld_h_n
port 1623 nsew signal input
flabel metal2 s 121848 996690 121900 996890 0 FreeSans 320 90 0 0 gpio4_5_analog_sel
port 1624 nsew signal input
flabel metal2 s 121497 996690 121549 996890 0 FreeSans 320 90 0 0 gpio4_5_dm[2]
port 1625 nsew signal input
flabel metal2 s 129166 996690 129218 996890 0 FreeSans 320 90 0 0 gpio4_5_dm[1]
port 1626 nsew signal input
flabel metal2 s 125770 996690 125822 996890 0 FreeSans 320 90 0 0 gpio4_5_dm[0]
port 1627 nsew signal input
flabel metal2 s 121119 996690 121171 996890 0 FreeSans 320 90 0 0 gpio4_5_hld_ovr
port 1628 nsew signal input
flabel metal2 s 120270 996690 120322 996890 0 FreeSans 320 90 0 0 gpio4_5_out
port 1629 nsew signal input
flabel metal2 s 119061 996690 119113 996890 0 FreeSans 320 90 0 0 gpio4_5_enable_vswitch_h
port 1630 nsew signal input
flabel metal2 s 118350 996690 118402 996890 0 FreeSans 320 90 0 0 gpio4_5_enable_vdda_h
port 1631 nsew signal input
flabel metal2 s 117102 996690 117154 996890 0 FreeSans 320 90 0 0 gpio4_5_vtrip_sel
port 1632 nsew signal input
flabel metal2 s 116782 996690 116834 996890 0 FreeSans 320 90 0 0 gpio4_5_ib_mode_sel
port 1633 nsew signal input
flabel metal2 s 116468 996690 116520 996890 0 FreeSans 320 90 0 0 gpio4_5_oe_n
port 1634 nsew signal input
flabel metal2 s 115878 996690 116002 996890 0 FreeSans 320 90 0 0 gpio4_5_in_h
port 1635 nsew signal input
flabel metal2 s 133254 996690 133306 996890 0 FreeSans 320 90 0 0 gpio4_5_zero
port 1636 nsew signal output
flabel metal2 s 133616 996690 133668 996890 0 FreeSans 320 90 0 0 gpio4_5_one
port 1637 nsew signal output
flabel metal2 s 108290 996690 108342 996890 0 FreeSans 320 90 0 0 gpio4_6_tie_lo_esd
port 1638 nsew signal output
flabel metal2 s 107990 996690 108042 996890 0 FreeSans 320 90 0 0 gpio4_6_in
port 1639 nsew signal output
flabel metal2 s 107688 996690 107740 996890 0 FreeSans 320 90 0 0 gpio4_6_tie_hi_esd
port 1640 nsew signal output
flabel metal2 s 107390 996690 107442 996890 0 FreeSans 320 90 0 0 gpio4_6_enable_vddio
port 1641 nsew signal input
flabel metal2 s 107090 996690 107142 996890 0 FreeSans 320 90 0 0 gpio4_6_slow
port 1642 nsew signal input
flabel metal2 s 106714 996690 106842 996890 0 FreeSans 320 90 0 0 gpio4_6_pad_a_esd_0_h
port 1643 nsew signal bidirectional
flabel metal2 s 105454 996690 105584 996890 0 FreeSans 320 90 0 0 gpio4_6_pad_a_esd_1_h
port 1644 nsew signal bidirectional
flabel metal2 s 104362 996690 104576 996890 0 FreeSans 320 90 0 0 gpio4_6_pad_a_noesd_h
port 1645 nsew signal bidirectional
flabel metal2 s 104058 996690 104110 996890 0 FreeSans 320 90 0 0 gpio4_6_analog_en
port 1646 nsew signal input
flabel metal2 s 101144 996690 101196 996890 0 FreeSans 320 90 0 0 gpio4_6_analog_pol
port 1647 nsew signal input
flabel metal2 s 100848 996690 100900 996890 0 FreeSans 320 90 0 0 gpio4_6_inp_dis
port 1648 nsew signal input
flabel metal2 s 99473 996690 99529 996890 0 FreeSans 320 90 0 0 gpio4_6_enable_inp_h
port 1649 nsew signal input
flabel metal2 s 98891 996690 98943 996890 0 FreeSans 320 90 0 0 gpio4_6_enable_h
port 1650 nsew signal input
flabel metal2 s 98162 996690 98214 996890 0 FreeSans 320 90 0 0 gpio4_6_hld_h_n
port 1651 nsew signal input
flabel metal2 s 97848 996690 97900 996890 0 FreeSans 320 90 0 0 gpio4_6_analog_sel
port 1652 nsew signal input
flabel metal2 s 97497 996690 97549 996890 0 FreeSans 320 90 0 0 gpio4_6_dm[2]
port 1653 nsew signal input
flabel metal2 s 105166 996690 105218 996890 0 FreeSans 320 90 0 0 gpio4_6_dm[1]
port 1654 nsew signal input
flabel metal2 s 101770 996690 101822 996890 0 FreeSans 320 90 0 0 gpio4_6_dm[0]
port 1655 nsew signal input
flabel metal2 s 97119 996690 97171 996890 0 FreeSans 320 90 0 0 gpio4_6_hld_ovr
port 1656 nsew signal input
flabel metal2 s 96270 996690 96322 996890 0 FreeSans 320 90 0 0 gpio4_6_out
port 1657 nsew signal input
flabel metal2 s 95061 996690 95113 996890 0 FreeSans 320 90 0 0 gpio4_6_enable_vswitch_h
port 1658 nsew signal input
flabel metal2 s 94350 996690 94402 996890 0 FreeSans 320 90 0 0 gpio4_6_enable_vdda_h
port 1659 nsew signal input
flabel metal2 s 93102 996690 93154 996890 0 FreeSans 320 90 0 0 gpio4_6_vtrip_sel
port 1660 nsew signal input
flabel metal2 s 92782 996690 92834 996890 0 FreeSans 320 90 0 0 gpio4_6_ib_mode_sel
port 1661 nsew signal input
flabel metal2 s 92468 996690 92520 996890 0 FreeSans 320 90 0 0 gpio4_6_oe_n
port 1662 nsew signal input
flabel metal2 s 91878 996690 92002 996890 0 FreeSans 320 90 0 0 gpio4_6_in_h
port 1663 nsew signal input
flabel metal2 s 109254 996690 109306 996890 0 FreeSans 320 90 0 0 gpio4_6_zero
port 1664 nsew signal output
flabel metal2 s 109616 996690 109668 996890 0 FreeSans 320 90 0 0 gpio4_6_one
port 1665 nsew signal output
flabel metal2 s 84290 996690 84342 996890 0 FreeSans 320 90 0 0 gpio4_7_tie_lo_esd
port 1666 nsew signal output
flabel metal2 s 83990 996690 84042 996890 0 FreeSans 320 90 0 0 gpio4_7_in
port 1667 nsew signal output
flabel metal2 s 83688 996690 83740 996890 0 FreeSans 320 90 0 0 gpio4_7_tie_hi_esd
port 1668 nsew signal output
flabel metal2 s 83390 996690 83442 996890 0 FreeSans 320 90 0 0 gpio4_7_enable_vddio
port 1669 nsew signal input
flabel metal2 s 83090 996690 83142 996890 0 FreeSans 320 90 0 0 gpio4_7_slow
port 1670 nsew signal input
flabel metal2 s 82714 996690 82842 996890 0 FreeSans 320 90 0 0 gpio4_7_pad_a_esd_0_h
port 1671 nsew signal bidirectional
flabel metal2 s 81454 996690 81584 996890 0 FreeSans 320 90 0 0 gpio4_7_pad_a_esd_1_h
port 1672 nsew signal bidirectional
flabel metal2 s 80362 996690 80576 996890 0 FreeSans 320 90 0 0 gpio4_7_pad_a_noesd_h
port 1673 nsew signal bidirectional
flabel metal2 s 80058 996690 80110 996890 0 FreeSans 320 90 0 0 gpio4_7_analog_en
port 1674 nsew signal input
flabel metal2 s 77144 996690 77196 996890 0 FreeSans 320 90 0 0 gpio4_7_analog_pol
port 1675 nsew signal input
flabel metal2 s 76848 996690 76900 996890 0 FreeSans 320 90 0 0 gpio4_7_inp_dis
port 1676 nsew signal input
flabel metal2 s 75473 996690 75529 996890 0 FreeSans 320 90 0 0 gpio4_7_enable_inp_h
port 1677 nsew signal input
flabel metal2 s 74891 996690 74943 996890 0 FreeSans 320 90 0 0 gpio4_7_enable_h
port 1678 nsew signal input
flabel metal2 s 74162 996690 74214 996890 0 FreeSans 320 90 0 0 gpio4_7_hld_h_n
port 1679 nsew signal input
flabel metal2 s 73848 996690 73900 996890 0 FreeSans 320 90 0 0 gpio4_7_analog_sel
port 1680 nsew signal input
flabel metal2 s 73497 996690 73549 996890 0 FreeSans 320 90 0 0 gpio4_7_dm[2]
port 1681 nsew signal input
flabel metal2 s 81166 996690 81218 996890 0 FreeSans 320 90 0 0 gpio4_7_dm[1]
port 1682 nsew signal input
flabel metal2 s 77770 996690 77822 996890 0 FreeSans 320 90 0 0 gpio4_7_dm[0]
port 1683 nsew signal input
flabel metal2 s 73119 996690 73171 996890 0 FreeSans 320 90 0 0 gpio4_7_hld_ovr
port 1684 nsew signal input
flabel metal2 s 72270 996690 72322 996890 0 FreeSans 320 90 0 0 gpio4_7_out
port 1685 nsew signal input
flabel metal2 s 71061 996690 71113 996890 0 FreeSans 320 90 0 0 gpio4_7_enable_vswitch_h
port 1686 nsew signal input
flabel metal2 s 70350 996690 70402 996890 0 FreeSans 320 90 0 0 gpio4_7_enable_vdda_h
port 1687 nsew signal input
flabel metal2 s 69102 996690 69154 996890 0 FreeSans 320 90 0 0 gpio4_7_vtrip_sel
port 1688 nsew signal input
flabel metal2 s 68782 996690 68834 996890 0 FreeSans 320 90 0 0 gpio4_7_ib_mode_sel
port 1689 nsew signal input
flabel metal2 s 68468 996690 68520 996890 0 FreeSans 320 90 0 0 gpio4_7_oe_n
port 1690 nsew signal input
flabel metal2 s 67878 996690 68002 996890 0 FreeSans 320 90 0 0 gpio4_7_in_h
port 1691 nsew signal input
flabel metal2 s 85254 996690 85306 996890 0 FreeSans 320 90 0 0 gpio4_7_zero
port 1692 nsew signal output
flabel metal2 s 85616 996690 85668 996890 0 FreeSans 320 90 0 0 gpio4_7_one
port 1693 nsew signal output
flabel metal3 s 40600 995154 40900 995214 0 FreeSans 320 0 0 0 muxsplit_nw_hld_vdda_h_n
port 1694 nsew signal input
flabel metal3 s 40600 994274 40900 994334 0 FreeSans 320 0 0 0 muxsplit_nw_enable_vdda_h
port 1695 nsew signal input
flabel metal3 s 40600 990652 40900 990712 0 FreeSans 320 0 0 0 muxsplit_nw_switch_aa_sl
port 1696 nsew signal input
flabel metal3 s 40600 990400 40900 990460 0 FreeSans 320 0 0 0 muxsplit_nw_switch_aa_s0
port 1697 nsew signal input
flabel metal3 s 40600 990148 40900 990208 0 FreeSans 320 0 0 0 muxsplit_nw_switch_bb_s0
port 1698 nsew signal input
flabel metal3 s 40600 989896 40900 989956 0 FreeSans 320 0 0 0 muxsplit_nw_switch_bb_sl
port 1699 nsew signal input
flabel metal3 s 40600 989644 40900 989704 0 FreeSans 320 0 0 0 muxsplit_nw_switch_bb_sr
port 1700 nsew signal input
flabel metal3 s 40600 989308 40900 989368 0 FreeSans 320 0 0 0 muxsplit_nw_switch_aa_sr
port 1701 nsew signal input
flabel metal3 s 40542 944602 40842 944672 0 FreeSans 320 0 0 0 gpio5_0_tie_lo_esd
port 1702 nsew signal output
flabel metal3 s 40538 944024 40838 944094 0 FreeSans 320 0 0 0 gpio5_0_in
port 1703 nsew signal output
flabel metal3 s 40542 944304 40842 944374 0 FreeSans 320 0 0 0 gpio5_0_tie_hi_esd
port 1704 nsew signal output
flabel metal3 s 40542 943712 40842 943782 0 FreeSans 320 0 0 0 gpio5_0_enable_vddio
port 1705 nsew signal input
flabel metal3 s 40542 943438 40842 943508 0 FreeSans 320 0 0 0 gpio5_0_slow
port 1706 nsew signal input
flabel metal3 s 40542 943090 40842 943218 0 FreeSans 320 0 0 0 gpio5_0_pad_a_esd_0_h
port 1707 nsew signal bidirectional
flabel metal3 s 40542 941658 40842 941788 0 FreeSans 320 0 0 0 gpio5_0_pad_a_esd_1_h
port 1708 nsew signal bidirectional
flabel metal3 s 40542 940564 40842 940778 0 FreeSans 320 0 0 0 gpio5_0_pad_a_noesd_h
port 1709 nsew signal bidirectional
flabel metal3 s 40542 939932 40842 940002 0 FreeSans 320 0 0 0 gpio5_0_analog_en
port 1710 nsew signal input
flabel metal3 s 40542 937172 40842 937242 0 FreeSans 320 0 0 0 gpio5_0_analog_pol
port 1711 nsew signal input
flabel metal3 s 40542 936592 40842 936662 0 FreeSans 320 0 0 0 gpio5_0_inp_dis
port 1712 nsew signal input
flabel metal3 s 40542 935426 40842 935496 0 FreeSans 320 0 0 0 gpio5_0_enable_inp_h
port 1713 nsew signal input
flabel metal3 s 40542 934970 40842 935040 0 FreeSans 320 0 0 0 gpio5_0_enable_h
port 1714 nsew signal input
flabel metal3 s 40542 934516 40842 934586 0 FreeSans 320 0 0 0 gpio5_0_hld_h_n
port 1715 nsew signal input
flabel metal3 s 40542 933898 40842 933968 0 FreeSans 320 0 0 0 gpio5_0_analog_sel
port 1716 nsew signal input
flabel metal3 s 40542 933454 40842 933524 0 FreeSans 320 0 0 0 gpio5_0_dm[2]
port 1717 nsew signal input
flabel metal3 s 40542 941128 40842 941198 0 FreeSans 320 0 0 0 gpio5_0_dm[1]
port 1718 nsew signal input
flabel metal3 s 40542 937720 40842 937790 0 FreeSans 320 0 0 0 gpio5_0_dm[0]
port 1719 nsew signal input
flabel metal3 s 40542 932970 40842 933040 0 FreeSans 320 0 0 0 gpio5_0_hld_ovr
port 1720 nsew signal input
flabel metal3 s 40542 932198 40842 932268 0 FreeSans 320 0 0 0 gpio5_0_out
port 1721 nsew signal input
flabel metal3 s 40542 930998 40842 931068 0 FreeSans 320 0 0 0 gpio5_0_enable_vswitch_h
port 1722 nsew signal input
flabel metal3 s 40542 930278 40842 930348 0 FreeSans 320 0 0 0 gpio5_0_enable_vdda_h
port 1723 nsew signal input
flabel metal3 s 40542 929416 40842 929486 0 FreeSans 320 0 0 0 gpio5_0_vtrip_sel
port 1724 nsew signal input
flabel metal3 s 40542 929072 40842 929142 0 FreeSans 320 0 0 0 gpio5_0_ib_mode_sel
port 1725 nsew signal input
flabel metal3 s 40542 928662 40842 928732 0 FreeSans 320 0 0 0 gpio5_0_oe_n
port 1726 nsew signal input
flabel metal3 s 40542 928080 40842 928204 0 FreeSans 320 0 0 0 gpio5_0_in_h
port 1727 nsew signal output
flabel metal3 s 40542 945802 40842 945872 0 FreeSans 320 0 0 0 gpio5_0_zero
port 1728 nsew signal output
flabel metal3 s 40542 946252 40842 946322 0 FreeSans 320 0 0 0 gpio5_0_one
port 1729 nsew signal output
flabel metal3 s 40542 923602 40842 923672 0 FreeSans 320 0 0 0 gpio5_1_tie_lo_esd
port 1730 nsew signal output
flabel metal3 s 40538 923024 40838 923094 0 FreeSans 320 0 0 0 gpio5_1_in
port 1731 nsew signal output
flabel metal3 s 40542 923304 40842 923374 0 FreeSans 320 0 0 0 gpio5_1_tie_hi_esd
port 1732 nsew signal output
flabel metal3 s 40542 922712 40842 922782 0 FreeSans 320 0 0 0 gpio5_1_enable_vddio
port 1733 nsew signal input
flabel metal3 s 40542 922438 40842 922508 0 FreeSans 320 0 0 0 gpio5_1_slow
port 1734 nsew signal input
flabel metal3 s 40542 922090 40842 922218 0 FreeSans 320 0 0 0 gpio5_1_pad_a_esd_0_h
port 1735 nsew signal bidirectional
flabel metal3 s 40542 920658 40842 920788 0 FreeSans 320 0 0 0 gpio5_1_pad_a_esd_1_h
port 1736 nsew signal bidirectional
flabel metal3 s 40542 919564 40842 919778 0 FreeSans 320 0 0 0 gpio5_1_pad_a_noesd_h
port 1737 nsew signal bidirectional
flabel metal3 s 40542 918932 40842 919002 0 FreeSans 320 0 0 0 gpio5_1_analog_en
port 1738 nsew signal input
flabel metal3 s 40542 916172 40842 916242 0 FreeSans 320 0 0 0 gpio5_1_analog_pol
port 1739 nsew signal input
flabel metal3 s 40542 915592 40842 915662 0 FreeSans 320 0 0 0 gpio5_1_inp_dis
port 1740 nsew signal input
flabel metal3 s 40542 914426 40842 914496 0 FreeSans 320 0 0 0 gpio5_1_enable_inp_h
port 1741 nsew signal input
flabel metal3 s 40542 913970 40842 914040 0 FreeSans 320 0 0 0 gpio5_1_enable_h
port 1742 nsew signal input
flabel metal3 s 40542 913516 40842 913586 0 FreeSans 320 0 0 0 gpio5_1_hld_h_n
port 1743 nsew signal input
flabel metal3 s 40542 912898 40842 912968 0 FreeSans 320 0 0 0 gpio5_1_analog_sel
port 1744 nsew signal input
flabel metal3 s 40542 912454 40842 912524 0 FreeSans 320 0 0 0 gpio5_1_dm[2]
port 1745 nsew signal input
flabel metal3 s 40542 920128 40842 920198 0 FreeSans 320 0 0 0 gpio5_1_dm[1]
port 1746 nsew signal input
flabel metal3 s 40542 916720 40842 916790 0 FreeSans 320 0 0 0 gpio5_1_dm[0]
port 1747 nsew signal input
flabel metal3 s 40542 911970 40842 912040 0 FreeSans 320 0 0 0 gpio5_1_hld_ovr
port 1748 nsew signal input
flabel metal3 s 40542 911198 40842 911268 0 FreeSans 320 0 0 0 gpio5_1_out
port 1749 nsew signal input
flabel metal3 s 40542 909998 40842 910068 0 FreeSans 320 0 0 0 gpio5_1_enable_vswitch_h
port 1750 nsew signal input
flabel metal3 s 40542 909278 40842 909348 0 FreeSans 320 0 0 0 gpio5_1_enable_vdda_h
port 1751 nsew signal input
flabel metal3 s 40542 908416 40842 908486 0 FreeSans 320 0 0 0 gpio5_1_vtrip_sel
port 1752 nsew signal input
flabel metal3 s 40542 908072 40842 908142 0 FreeSans 320 0 0 0 gpio5_1_ib_mode_sel
port 1753 nsew signal input
flabel metal3 s 40542 907662 40842 907732 0 FreeSans 320 0 0 0 gpio5_1_oe_n
port 1754 nsew signal input
flabel metal3 s 40542 907080 40842 907204 0 FreeSans 320 0 0 0 gpio5_1_in_h
port 1755 nsew signal output
flabel metal3 s 40542 924802 40842 924872 0 FreeSans 320 0 0 0 gpio5_1_zero
port 1756 nsew signal output
flabel metal3 s 40542 925252 40842 925322 0 FreeSans 320 0 0 0 gpio5_1_one
port 1757 nsew signal output
flabel metal3 s 40542 902602 40842 902672 0 FreeSans 320 0 0 0 gpio5_2_tie_lo_esd
port 1758 nsew signal output
flabel metal3 s 40538 902024 40838 902094 0 FreeSans 320 0 0 0 gpio5_2_in
port 1759 nsew signal output
flabel metal3 s 40542 902304 40842 902374 0 FreeSans 320 0 0 0 gpio5_2_tie_hi_esd
port 1760 nsew signal output
flabel metal3 s 40542 901712 40842 901782 0 FreeSans 320 0 0 0 gpio5_2_enable_vddio
port 1761 nsew signal input
flabel metal3 s 40542 901438 40842 901508 0 FreeSans 320 0 0 0 gpio5_2_slow
port 1762 nsew signal input
flabel metal3 s 40542 901090 40842 901218 0 FreeSans 320 0 0 0 gpio5_2_pad_a_esd_0_h
port 1763 nsew signal bidirectional
flabel metal3 s 40542 899658 40842 899788 0 FreeSans 320 0 0 0 gpio5_2_pad_a_esd_1_h
port 1764 nsew signal bidirectional
flabel metal3 s 40542 898564 40842 898778 0 FreeSans 320 0 0 0 gpio5_2_pad_a_noesd_h
port 1765 nsew signal bidirectional
flabel metal3 s 40542 897932 40842 898002 0 FreeSans 320 0 0 0 gpio5_2_analog_en
port 1766 nsew signal input
flabel metal3 s 40542 895172 40842 895242 0 FreeSans 320 0 0 0 gpio5_2_analog_pol
port 1767 nsew signal input
flabel metal3 s 40542 894592 40842 894662 0 FreeSans 320 0 0 0 gpio5_2_inp_dis
port 1768 nsew signal input
flabel metal3 s 40542 893426 40842 893496 0 FreeSans 320 0 0 0 gpio5_2_enable_inp_h
port 1769 nsew signal input
flabel metal3 s 40542 892970 40842 893040 0 FreeSans 320 0 0 0 gpio5_2_enable_h
port 1770 nsew signal input
flabel metal3 s 40542 892516 40842 892586 0 FreeSans 320 0 0 0 gpio5_2_hld_h_n
port 1771 nsew signal input
flabel metal3 s 40542 891898 40842 891968 0 FreeSans 320 0 0 0 gpio5_2_analog_sel
port 1772 nsew signal input
flabel metal3 s 40542 891454 40842 891524 0 FreeSans 320 0 0 0 gpio5_2_dm[2]
port 1773 nsew signal input
flabel metal3 s 40542 899128 40842 899198 0 FreeSans 320 0 0 0 gpio5_2_dm[1]
port 1774 nsew signal input
flabel metal3 s 40542 895720 40842 895790 0 FreeSans 320 0 0 0 gpio5_2_dm[0]
port 1775 nsew signal input
flabel metal3 s 40542 890970 40842 891040 0 FreeSans 320 0 0 0 gpio5_2_hld_ovr
port 1776 nsew signal input
flabel metal3 s 40542 890198 40842 890268 0 FreeSans 320 0 0 0 gpio5_2_out
port 1777 nsew signal input
flabel metal3 s 40542 888998 40842 889068 0 FreeSans 320 0 0 0 gpio5_2_enable_vswitch_h
port 1778 nsew signal input
flabel metal3 s 40542 888278 40842 888348 0 FreeSans 320 0 0 0 gpio5_2_enable_vdda_h
port 1779 nsew signal input
flabel metal3 s 40542 887416 40842 887486 0 FreeSans 320 0 0 0 gpio5_2_vtrip_sel
port 1780 nsew signal input
flabel metal3 s 40542 887072 40842 887142 0 FreeSans 320 0 0 0 gpio5_2_ib_mode_sel
port 1781 nsew signal input
flabel metal3 s 40542 886662 40842 886732 0 FreeSans 320 0 0 0 gpio5_2_oe_n
port 1782 nsew signal input
flabel metal3 s 40542 886080 40842 886204 0 FreeSans 320 0 0 0 gpio5_2_in_h
port 1783 nsew signal output
flabel metal3 s 40542 903802 40842 903872 0 FreeSans 320 0 0 0 gpio5_2_zero
port 1784 nsew signal output
flabel metal3 s 40542 904252 40842 904322 0 FreeSans 320 0 0 0 gpio5_2_one
port 1785 nsew signal output
flabel metal3 s 40542 881602 40842 881672 0 FreeSans 320 0 0 0 gpio5_3_tie_lo_esd
port 1786 nsew signal output
flabel metal3 s 40538 881024 40838 881094 0 FreeSans 320 0 0 0 gpio5_3_in
port 1787 nsew signal output
flabel metal3 s 40542 881304 40842 881374 0 FreeSans 320 0 0 0 gpio5_3_tie_hi_esd
port 1788 nsew signal output
flabel metal3 s 40542 880712 40842 880782 0 FreeSans 320 0 0 0 gpio5_3_enable_vddio
port 1789 nsew signal input
flabel metal3 s 40542 880438 40842 880508 0 FreeSans 320 0 0 0 gpio5_3_slow
port 1790 nsew signal input
flabel metal3 s 40542 880090 40842 880218 0 FreeSans 320 0 0 0 gpio5_3_pad_a_esd_0_h
port 1791 nsew signal bidirectional
flabel metal3 s 40542 878658 40842 878788 0 FreeSans 320 0 0 0 gpio5_3_pad_a_esd_1_h
port 1792 nsew signal bidirectional
flabel metal3 s 40542 877564 40842 877778 0 FreeSans 320 0 0 0 gpio5_3_pad_a_noesd_h
port 1793 nsew signal bidirectional
flabel metal3 s 40542 876932 40842 877002 0 FreeSans 320 0 0 0 gpio5_3_analog_en
port 1794 nsew signal input
flabel metal3 s 40542 874172 40842 874242 0 FreeSans 320 0 0 0 gpio5_3_analog_pol
port 1795 nsew signal input
flabel metal3 s 40542 873592 40842 873662 0 FreeSans 320 0 0 0 gpio5_3_inp_dis
port 1796 nsew signal input
flabel metal3 s 40542 872426 40842 872496 0 FreeSans 320 0 0 0 gpio5_3_enable_inp_h
port 1797 nsew signal input
flabel metal3 s 40542 871970 40842 872040 0 FreeSans 320 0 0 0 gpio5_3_enable_h
port 1798 nsew signal input
flabel metal3 s 40542 871516 40842 871586 0 FreeSans 320 0 0 0 gpio5_3_hld_h_n
port 1799 nsew signal input
flabel metal3 s 40542 870898 40842 870968 0 FreeSans 320 0 0 0 gpio5_3_analog_sel
port 1800 nsew signal input
flabel metal3 s 40542 870454 40842 870524 0 FreeSans 320 0 0 0 gpio5_3_dm[2]
port 1801 nsew signal input
flabel metal3 s 40542 878128 40842 878198 0 FreeSans 320 0 0 0 gpio5_3_dm[1]
port 1802 nsew signal input
flabel metal3 s 40542 874720 40842 874790 0 FreeSans 320 0 0 0 gpio5_3_dm[0]
port 1803 nsew signal input
flabel metal3 s 40542 869970 40842 870040 0 FreeSans 320 0 0 0 gpio5_3_hld_ovr
port 1804 nsew signal input
flabel metal3 s 40542 869198 40842 869268 0 FreeSans 320 0 0 0 gpio5_3_out
port 1805 nsew signal input
flabel metal3 s 40542 867998 40842 868068 0 FreeSans 320 0 0 0 gpio5_3_enable_vswitch_h
port 1806 nsew signal input
flabel metal3 s 40542 867278 40842 867348 0 FreeSans 320 0 0 0 gpio5_3_enable_vdda_h
port 1807 nsew signal input
flabel metal3 s 40542 866416 40842 866486 0 FreeSans 320 0 0 0 gpio5_3_vtrip_sel
port 1808 nsew signal input
flabel metal3 s 40542 866072 40842 866142 0 FreeSans 320 0 0 0 gpio5_3_ib_mode_sel
port 1809 nsew signal input
flabel metal3 s 40542 865662 40842 865732 0 FreeSans 320 0 0 0 gpio5_3_oe_n
port 1810 nsew signal input
flabel metal3 s 40542 865080 40842 865204 0 FreeSans 320 0 0 0 gpio5_3_in_h
port 1811 nsew signal output
flabel metal3 s 40542 882802 40842 882872 0 FreeSans 320 0 0 0 gpio5_3_zero
port 1812 nsew signal output
flabel metal3 s 40542 883252 40842 883322 0 FreeSans 320 0 0 0 gpio5_3_one
port 1813 nsew signal output
flabel metal3 s 40542 840602 40842 840672 0 FreeSans 320 0 0 0 gpio5_4_tie_lo_esd
port 1814 nsew signal output
flabel metal3 s 40538 840024 40838 840094 0 FreeSans 320 0 0 0 gpio5_4_in
port 1815 nsew signal output
flabel metal3 s 40542 840304 40842 840374 0 FreeSans 320 0 0 0 gpio5_4_tie_hi_esd
port 1816 nsew signal output
flabel metal3 s 40542 839712 40842 839782 0 FreeSans 320 0 0 0 gpio5_4_enable_vddio
port 1817 nsew signal input
flabel metal3 s 40542 839438 40842 839508 0 FreeSans 320 0 0 0 gpio5_4_slow
port 1818 nsew signal input
flabel metal3 s 40542 839090 40842 839218 0 FreeSans 320 0 0 0 gpio5_4_pad_a_esd_0_h
port 1819 nsew signal bidirectional
flabel metal3 s 40542 837658 40842 837788 0 FreeSans 320 0 0 0 gpio5_4_pad_a_esd_1_h
port 1820 nsew signal bidirectional
flabel metal3 s 40542 836564 40842 836778 0 FreeSans 320 0 0 0 gpio5_4_pad_a_noesd_h
port 1821 nsew signal bidirectional
flabel metal3 s 40542 835932 40842 836002 0 FreeSans 320 0 0 0 gpio5_4_analog_en
port 1822 nsew signal input
flabel metal3 s 40542 833172 40842 833242 0 FreeSans 320 0 0 0 gpio5_4_analog_pol
port 1823 nsew signal input
flabel metal3 s 40542 832592 40842 832662 0 FreeSans 320 0 0 0 gpio5_4_inp_dis
port 1824 nsew signal input
flabel metal3 s 40542 831426 40842 831496 0 FreeSans 320 0 0 0 gpio5_4_enable_inp_h
port 1825 nsew signal input
flabel metal3 s 40542 830970 40842 831040 0 FreeSans 320 0 0 0 gpio5_4_enable_h
port 1826 nsew signal input
flabel metal3 s 40542 830516 40842 830586 0 FreeSans 320 0 0 0 gpio5_4_hld_h_n
port 1827 nsew signal input
flabel metal3 s 40542 829898 40842 829968 0 FreeSans 320 0 0 0 gpio5_4_analog_sel
port 1828 nsew signal input
flabel metal3 s 40542 829454 40842 829524 0 FreeSans 320 0 0 0 gpio5_4_dm[2]
port 1829 nsew signal input
flabel metal3 s 40542 837128 40842 837198 0 FreeSans 320 0 0 0 gpio5_4_dm[1]
port 1830 nsew signal input
flabel metal3 s 40542 833720 40842 833790 0 FreeSans 320 0 0 0 gpio5_4_dm[0]
port 1831 nsew signal input
flabel metal3 s 40542 828970 40842 829040 0 FreeSans 320 0 0 0 gpio5_4_hld_ovr
port 1832 nsew signal input
flabel metal3 s 40542 828198 40842 828268 0 FreeSans 320 0 0 0 gpio5_4_out
port 1833 nsew signal input
flabel metal3 s 40542 826998 40842 827068 0 FreeSans 320 0 0 0 gpio5_4_enable_vswitch_h
port 1834 nsew signal input
flabel metal3 s 40542 826278 40842 826348 0 FreeSans 320 0 0 0 gpio5_4_enable_vdda_h
port 1835 nsew signal input
flabel metal3 s 40542 825416 40842 825486 0 FreeSans 320 0 0 0 gpio5_4_vtrip_sel
port 1836 nsew signal input
flabel metal3 s 40542 825072 40842 825142 0 FreeSans 320 0 0 0 gpio5_4_ib_mode_sel
port 1837 nsew signal input
flabel metal3 s 40542 824662 40842 824732 0 FreeSans 320 0 0 0 gpio5_4_oe_n
port 1838 nsew signal input
flabel metal3 s 40542 824080 40842 824204 0 FreeSans 320 0 0 0 gpio5_4_in_h
port 1839 nsew signal output
flabel metal3 s 40542 841802 40842 841872 0 FreeSans 320 0 0 0 gpio5_4_zero
port 1840 nsew signal output
flabel metal3 s 40542 842252 40842 842322 0 FreeSans 320 0 0 0 gpio5_4_one
port 1841 nsew signal output
flabel metal3 s 40542 819602 40842 819672 0 FreeSans 320 0 0 0 gpio5_5_tie_lo_esd
port 1842 nsew signal output
flabel metal3 s 40538 819024 40838 819094 0 FreeSans 320 0 0 0 gpio5_5_in
port 1843 nsew signal output
flabel metal3 s 40542 819304 40842 819374 0 FreeSans 320 0 0 0 gpio5_5_tie_hi_esd
port 1844 nsew signal output
flabel metal3 s 40542 818712 40842 818782 0 FreeSans 320 0 0 0 gpio5_5_enable_vddio
port 1845 nsew signal input
flabel metal3 s 40542 818438 40842 818508 0 FreeSans 320 0 0 0 gpio5_5_slow
port 1846 nsew signal input
flabel metal3 s 40542 818090 40842 818218 0 FreeSans 320 0 0 0 gpio5_5_pad_a_esd_0_h
port 1847 nsew signal bidirectional
flabel metal3 s 40542 816658 40842 816788 0 FreeSans 320 0 0 0 gpio5_5_pad_a_esd_1_h
port 1848 nsew signal bidirectional
flabel metal3 s 40542 815564 40842 815778 0 FreeSans 320 0 0 0 gpio5_5_pad_a_noesd_h
port 1849 nsew signal bidirectional
flabel metal3 s 40542 814932 40842 815002 0 FreeSans 320 0 0 0 gpio5_5_analog_en
port 1850 nsew signal input
flabel metal3 s 40542 812172 40842 812242 0 FreeSans 320 0 0 0 gpio5_5_analog_pol
port 1851 nsew signal input
flabel metal3 s 40542 811592 40842 811662 0 FreeSans 320 0 0 0 gpio5_5_inp_dis
port 1852 nsew signal input
flabel metal3 s 40542 810426 40842 810496 0 FreeSans 320 0 0 0 gpio5_5_enable_inp_h
port 1853 nsew signal input
flabel metal3 s 40542 809970 40842 810040 0 FreeSans 320 0 0 0 gpio5_5_enable_h
port 1854 nsew signal input
flabel metal3 s 40542 809516 40842 809586 0 FreeSans 320 0 0 0 gpio5_5_hld_h_n
port 1855 nsew signal input
flabel metal3 s 40542 808898 40842 808968 0 FreeSans 320 0 0 0 gpio5_5_analog_sel
port 1856 nsew signal input
flabel metal3 s 40542 808454 40842 808524 0 FreeSans 320 0 0 0 gpio5_5_dm[2]
port 1857 nsew signal input
flabel metal3 s 40542 816128 40842 816198 0 FreeSans 320 0 0 0 gpio5_5_dm[1]
port 1858 nsew signal input
flabel metal3 s 40542 812720 40842 812790 0 FreeSans 320 0 0 0 gpio5_5_dm[0]
port 1859 nsew signal input
flabel metal3 s 40542 807970 40842 808040 0 FreeSans 320 0 0 0 gpio5_5_hld_ovr
port 1860 nsew signal input
flabel metal3 s 40542 807198 40842 807268 0 FreeSans 320 0 0 0 gpio5_5_out
port 1861 nsew signal input
flabel metal3 s 40542 805998 40842 806068 0 FreeSans 320 0 0 0 gpio5_5_enable_vswitch_h
port 1862 nsew signal input
flabel metal3 s 40542 805278 40842 805348 0 FreeSans 320 0 0 0 gpio5_5_enable_vdda_h
port 1863 nsew signal input
flabel metal3 s 40542 804416 40842 804486 0 FreeSans 320 0 0 0 gpio5_5_vtrip_sel
port 1864 nsew signal input
flabel metal3 s 40542 804072 40842 804142 0 FreeSans 320 0 0 0 gpio5_5_ib_mode_sel
port 1865 nsew signal input
flabel metal3 s 40542 803662 40842 803732 0 FreeSans 320 0 0 0 gpio5_5_oe_n
port 1866 nsew signal input
flabel metal3 s 40542 803080 40842 803204 0 FreeSans 320 0 0 0 gpio5_5_in_h
port 1867 nsew signal output
flabel metal3 s 40542 820802 40842 820872 0 FreeSans 320 0 0 0 gpio5_5_zero
port 1868 nsew signal output
flabel metal3 s 40542 821252 40842 821322 0 FreeSans 320 0 0 0 gpio5_5_one
port 1869 nsew signal output
flabel metal3 s 40542 798602 40842 798672 0 FreeSans 320 0 0 0 gpio5_6_tie_lo_esd
port 1870 nsew signal output
flabel metal3 s 40538 798024 40838 798094 0 FreeSans 320 0 0 0 gpio5_6_in
port 1871 nsew signal output
flabel metal3 s 40542 798304 40842 798374 0 FreeSans 320 0 0 0 gpio5_6_tie_hi_esd
port 1872 nsew signal output
flabel metal3 s 40542 797712 40842 797782 0 FreeSans 320 0 0 0 gpio5_6_enable_vddio
port 1873 nsew signal input
flabel metal3 s 40542 797438 40842 797508 0 FreeSans 320 0 0 0 gpio5_6_slow
port 1874 nsew signal input
flabel metal3 s 40542 797090 40842 797218 0 FreeSans 320 0 0 0 gpio5_6_pad_a_esd_0_h
port 1875 nsew signal bidirectional
flabel metal3 s 40542 795658 40842 795788 0 FreeSans 320 0 0 0 gpio5_6_pad_a_esd_1_h
port 1876 nsew signal bidirectional
flabel metal3 s 40542 794564 40842 794778 0 FreeSans 320 0 0 0 gpio5_6_pad_a_noesd_h
port 1877 nsew signal bidirectional
flabel metal3 s 40542 793932 40842 794002 0 FreeSans 320 0 0 0 gpio5_6_analog_en
port 1878 nsew signal input
flabel metal3 s 40542 791172 40842 791242 0 FreeSans 320 0 0 0 gpio5_6_analog_pol
port 1879 nsew signal input
flabel metal3 s 40542 790592 40842 790662 0 FreeSans 320 0 0 0 gpio5_6_inp_dis
port 1880 nsew signal input
flabel metal3 s 40542 789426 40842 789496 0 FreeSans 320 0 0 0 gpio5_6_enable_inp_h
port 1881 nsew signal input
flabel metal3 s 40542 788970 40842 789040 0 FreeSans 320 0 0 0 gpio5_6_enable_h
port 1882 nsew signal input
flabel metal3 s 40542 788516 40842 788586 0 FreeSans 320 0 0 0 gpio5_6_hld_h_n
port 1883 nsew signal input
flabel metal3 s 40542 787898 40842 787968 0 FreeSans 320 0 0 0 gpio5_6_analog_sel
port 1884 nsew signal input
flabel metal3 s 40542 787454 40842 787524 0 FreeSans 320 0 0 0 gpio5_6_dm[2]
port 1885 nsew signal input
flabel metal3 s 40542 795128 40842 795198 0 FreeSans 320 0 0 0 gpio5_6_dm[1]
port 1886 nsew signal input
flabel metal3 s 40542 791720 40842 791790 0 FreeSans 320 0 0 0 gpio5_6_dm[0]
port 1887 nsew signal input
flabel metal3 s 40542 786970 40842 787040 0 FreeSans 320 0 0 0 gpio5_6_hld_ovr
port 1888 nsew signal input
flabel metal3 s 40542 786198 40842 786268 0 FreeSans 320 0 0 0 gpio5_6_out
port 1889 nsew signal input
flabel metal3 s 40542 784998 40842 785068 0 FreeSans 320 0 0 0 gpio5_6_enable_vswitch_h
port 1890 nsew signal input
flabel metal3 s 40542 784278 40842 784348 0 FreeSans 320 0 0 0 gpio5_6_enable_vdda_h
port 1891 nsew signal input
flabel metal3 s 40542 783416 40842 783486 0 FreeSans 320 0 0 0 gpio5_6_vtrip_sel
port 1892 nsew signal input
flabel metal3 s 40542 783072 40842 783142 0 FreeSans 320 0 0 0 gpio5_6_ib_mode_sel
port 1893 nsew signal input
flabel metal3 s 40542 782662 40842 782732 0 FreeSans 320 0 0 0 gpio5_6_oe_n
port 1894 nsew signal input
flabel metal3 s 40542 782080 40842 782204 0 FreeSans 320 0 0 0 gpio5_6_in_h
port 1895 nsew signal output
flabel metal3 s 40542 799802 40842 799872 0 FreeSans 320 0 0 0 gpio5_6_zero
port 1896 nsew signal output
flabel metal3 s 40542 800252 40842 800322 0 FreeSans 320 0 0 0 gpio5_6_one
port 1897 nsew signal output
flabel metal3 s 40542 777602 40842 777672 0 FreeSans 320 0 0 0 gpio5_7_tie_lo_esd
port 1898 nsew signal output
flabel metal3 s 40538 777024 40838 777094 0 FreeSans 320 0 0 0 gpio5_7_in
port 1899 nsew signal output
flabel metal3 s 40542 777304 40842 777374 0 FreeSans 320 0 0 0 gpio5_7_tie_hi_esd
port 1900 nsew signal output
flabel metal3 s 40542 776712 40842 776782 0 FreeSans 320 0 0 0 gpio5_7_enable_vddio
port 1901 nsew signal input
flabel metal3 s 40542 776438 40842 776508 0 FreeSans 320 0 0 0 gpio5_7_slow
port 1902 nsew signal input
flabel metal3 s 40542 776090 40842 776218 0 FreeSans 320 0 0 0 gpio5_7_pad_a_esd_0_h
port 1903 nsew signal bidirectional
flabel metal3 s 40542 774658 40842 774788 0 FreeSans 320 0 0 0 gpio5_7_pad_a_esd_1_h
port 1904 nsew signal bidirectional
flabel metal3 s 40542 773564 40842 773778 0 FreeSans 320 0 0 0 gpio5_7_pad_a_noesd_h
port 1905 nsew signal bidirectional
flabel metal3 s 40542 772932 40842 773002 0 FreeSans 320 0 0 0 gpio5_7_analog_en
port 1906 nsew signal input
flabel metal3 s 40542 770172 40842 770242 0 FreeSans 320 0 0 0 gpio5_7_analog_pol
port 1907 nsew signal input
flabel metal3 s 40542 769592 40842 769662 0 FreeSans 320 0 0 0 gpio5_7_inp_dis
port 1908 nsew signal input
flabel metal3 s 40542 768426 40842 768496 0 FreeSans 320 0 0 0 gpio5_7_enable_inp_h
port 1909 nsew signal input
flabel metal3 s 40542 767970 40842 768040 0 FreeSans 320 0 0 0 gpio5_7_enable_h
port 1910 nsew signal input
flabel metal3 s 40542 767516 40842 767586 0 FreeSans 320 0 0 0 gpio5_7_hld_h_n
port 1911 nsew signal input
flabel metal3 s 40542 766898 40842 766968 0 FreeSans 320 0 0 0 gpio5_7_analog_sel
port 1912 nsew signal input
flabel metal3 s 40542 766454 40842 766524 0 FreeSans 320 0 0 0 gpio5_7_dm[2]
port 1913 nsew signal input
flabel metal3 s 40542 774128 40842 774198 0 FreeSans 320 0 0 0 gpio5_7_dm[1]
port 1914 nsew signal input
flabel metal3 s 40542 770720 40842 770790 0 FreeSans 320 0 0 0 gpio5_7_dm[0]
port 1915 nsew signal input
flabel metal3 s 40542 765970 40842 766040 0 FreeSans 320 0 0 0 gpio5_7_hld_ovr
port 1916 nsew signal input
flabel metal3 s 40542 765198 40842 765268 0 FreeSans 320 0 0 0 gpio5_7_out
port 1917 nsew signal input
flabel metal3 s 40542 763998 40842 764068 0 FreeSans 320 0 0 0 gpio5_7_enable_vswitch_h
port 1918 nsew signal input
flabel metal3 s 40542 763278 40842 763348 0 FreeSans 320 0 0 0 gpio5_7_enable_vdda_h
port 1919 nsew signal input
flabel metal3 s 40542 762416 40842 762486 0 FreeSans 320 0 0 0 gpio5_7_vtrip_sel
port 1920 nsew signal input
flabel metal3 s 40542 762072 40842 762142 0 FreeSans 320 0 0 0 gpio5_7_ib_mode_sel
port 1921 nsew signal input
flabel metal3 s 40542 761662 40842 761732 0 FreeSans 320 0 0 0 gpio5_7_oe_n
port 1922 nsew signal input
flabel metal3 s 40542 761080 40842 761204 0 FreeSans 320 0 0 0 gpio5_7_in_h
port 1923 nsew signal output
flabel metal3 s 40542 778802 40842 778872 0 FreeSans 320 0 0 0 gpio5_7_zero
port 1924 nsew signal output
flabel metal3 s 40542 779252 40842 779322 0 FreeSans 320 0 0 0 gpio5_7_one
port 1925 nsew signal output
flabel metal3 s 40300 670995 40600 671061 0 FreeSans 320 0 0 0 gpio6_0_tie_hi_esd
port 1926 nsew signal output
flabel metal3 s 40300 666679 40600 666745 0 FreeSans 320 0 0 0 gpio6_0_dm[2]
port 1927 nsew signal input
flabel metal3 s 40300 670655 40600 670721 0 FreeSans 320 0 0 0 gpio6_0_dm[1]
port 1928 nsew signal input
flabel metal3 s 40300 670825 40600 670891 0 FreeSans 320 0 0 0 gpio6_0_dm[0]
port 1929 nsew signal input
flabel metal3 s 40300 670028 40600 670094 0 FreeSans 320 0 0 0 gpio6_0_slow
port 1930 nsew signal input
flabel metal3 s 40300 669889 40600 669955 0 FreeSans 320 0 0 0 gpio6_0_oe_n
port 1931 nsew signal input
flabel metal3 s 40300 668058 40600 668178 0 FreeSans 320 0 0 0 gpio6_0_tie_lo_esd
port 1932 nsew signal output
flabel metal3 s 40300 666509 40600 666575 0 FreeSans 320 0 0 0 gpio6_0_inp_dis
port 1933 nsew signal input
flabel metal3 s 40300 664169 40600 664243 0 FreeSans 320 0 0 0 gpio6_0_enable_vddio
port 1934 nsew signal input
flabel metal3 s 40300 662533 40600 662599 0 FreeSans 320 0 0 0 gpio6_0_vtrip_sel
port 1935 nsew signal input
flabel metal3 s 40300 658387 40600 658453 0 FreeSans 320 0 0 0 gpio6_0_ib_mode_sel[1]
port 1936 nsew signal input
flabel metal3 s 40300 662363 40600 662429 0 FreeSans 320 0 0 0 gpio6_0_ib_mode_sel[0]
port 1937 nsew signal input
flabel metal3 s 40300 659825 40600 659891 0 FreeSans 320 0 0 0 gpio6_0_out
port 1938 nsew signal input
flabel metal3 s 40300 654241 40600 654307 0 FreeSans 320 0 0 0 gpio6_0_slew_ctl[1]
port 1939 nsew signal input
flabel metal3 s 40300 658217 40600 658283 0 FreeSans 320 0 0 0 gpio6_0_slew_ctl[0]
port 1940 nsew signal input
flabel metal3 s 40300 658047 40600 658113 0 FreeSans 320 0 0 0 gpio6_0_analog_pol
port 1941 nsew signal input
flabel metal3 s 40300 655331 40600 655397 0 FreeSans 320 0 0 0 gpio6_0_analog_sel
port 1942 nsew signal input
flabel metal3 s 40300 654071 40600 654137 0 FreeSans 320 0 0 0 gpio6_0_hys_trim
port 1943 nsew signal input
flabel metal3 s 40300 653807 40600 653873 0 FreeSans 320 0 0 0 gpio6_0_vinref
port 1944 nsew signal input
flabel metal3 s 40300 650471 40600 650537 0 FreeSans 320 0 0 0 gpio6_0_hld_ovr
port 1945 nsew signal input
flabel metal3 s 40300 649876 40600 649942 0 FreeSans 320 0 0 0 gpio6_0_in_h
port 1946 nsew signal output
flabel metal3 s 40300 649427 40600 649493 0 FreeSans 320 0 0 0 gpio6_0_enable_h
port 1947 nsew signal input
flabel metal3 s 40300 649076 40600 649142 0 FreeSans 320 0 0 0 gpio6_0_in
port 1948 nsew signal output
flabel metal3 s 40300 648927 40600 648993 0 FreeSans 320 0 0 0 gpio6_0_hld_h_n
port 1949 nsew signal input
flabel metal3 s 40300 646754 40600 646820 0 FreeSans 320 0 0 0 gpio6_0_enable_vdda_h
port 1950 nsew signal input
flabel metal3 s 40300 646623 40600 646689 0 FreeSans 320 0 0 0 gpio6_0_analog_en
port 1951 nsew signal input
flabel metal3 s 40300 646422 40600 646488 0 FreeSans 320 0 0 0 gpio6_0_enable_inp_h
port 1952 nsew signal input
flabel metal3 s 40300 646153 40600 646273 0 FreeSans 320 0 0 0 gpio6_0_enable_vswitch_h
port 1953 nsew signal input
flabel metal3 s 40300 645577 40600 645697 0 FreeSans 320 0 0 0 gpio6_0_pad_a_noesd_h
port 1954 nsew signal bidirectional
flabel metal3 s 40300 645321 40600 645440 0 FreeSans 320 0 0 0 gpio6_0_pad_a_esd_0_h
port 1955 nsew signal bidirectional
flabel metal3 s 40300 645066 40600 645186 0 FreeSans 320 0 0 0 gpio6_0_pad_a_esd_1_h
port 1956 nsew signal bidirectional
flabel metal3 s 40300 674802 40600 674872 0 FreeSans 320 0 0 0 gpio6_0_zero
port 1957 nsew signal output
flabel metal3 s 40300 675252 40600 675322 0 FreeSans 320 0 0 0 gpio6_0_one
port 1958 nsew signal output
flabel metal3 s 40300 637995 40600 638061 0 FreeSans 320 0 0 0 gpio6_1_tie_hi_esd
port 1959 nsew signal output
flabel metal3 s 40300 633679 40600 633745 0 FreeSans 320 0 0 0 gpio6_1_dm[2]
port 1960 nsew signal input
flabel metal3 s 40300 637655 40600 637721 0 FreeSans 320 0 0 0 gpio6_1_dm[1]
port 1961 nsew signal input
flabel metal3 s 40300 637825 40600 637891 0 FreeSans 320 0 0 0 gpio6_1_dm[0]
port 1962 nsew signal input
flabel metal3 s 40300 637028 40600 637094 0 FreeSans 320 0 0 0 gpio6_1_slow
port 1963 nsew signal input
flabel metal3 s 40300 636889 40600 636955 0 FreeSans 320 0 0 0 gpio6_1_oe_n
port 1964 nsew signal input
flabel metal3 s 40300 635058 40600 635178 0 FreeSans 320 0 0 0 gpio6_1_tie_lo_esd
port 1965 nsew signal output
flabel metal3 s 40300 633509 40600 633575 0 FreeSans 320 0 0 0 gpio6_1_inp_dis
port 1966 nsew signal input
flabel metal3 s 40300 631169 40600 631243 0 FreeSans 320 0 0 0 gpio6_1_enable_vddio
port 1967 nsew signal input
flabel metal3 s 40300 629533 40600 629599 0 FreeSans 320 0 0 0 gpio6_1_vtrip_sel
port 1968 nsew signal input
flabel metal3 s 40300 625387 40600 625453 0 FreeSans 320 0 0 0 gpio6_1_ib_mode_sel[1]
port 1969 nsew signal input
flabel metal3 s 40300 629363 40600 629429 0 FreeSans 320 0 0 0 gpio6_1_ib_mode_sel[0]
port 1970 nsew signal input
flabel metal3 s 40300 626825 40600 626891 0 FreeSans 320 0 0 0 gpio6_1_out
port 1971 nsew signal input
flabel metal3 s 40300 621241 40600 621307 0 FreeSans 320 0 0 0 gpio6_1_slew_ctl[1]
port 1972 nsew signal input
flabel metal3 s 40300 625217 40600 625283 0 FreeSans 320 0 0 0 gpio6_1_slew_ctl[0]
port 1973 nsew signal input
flabel metal3 s 40300 625047 40600 625113 0 FreeSans 320 0 0 0 gpio6_1_analog_pol
port 1974 nsew signal input
flabel metal3 s 40300 622331 40600 622397 0 FreeSans 320 0 0 0 gpio6_1_analog_sel
port 1975 nsew signal input
flabel metal3 s 40300 621071 40600 621137 0 FreeSans 320 0 0 0 gpio6_1_hys_trim
port 1976 nsew signal input
flabel metal3 s 40300 620807 40600 620873 0 FreeSans 320 0 0 0 gpio6_1_vinref
port 1977 nsew signal input
flabel metal3 s 40300 617471 40600 617537 0 FreeSans 320 0 0 0 gpio6_1_hld_ovr
port 1978 nsew signal input
flabel metal3 s 40300 616876 40600 616942 0 FreeSans 320 0 0 0 gpio6_1_in_h
port 1979 nsew signal output
flabel metal3 s 40300 616427 40600 616493 0 FreeSans 320 0 0 0 gpio6_1_enable_h
port 1980 nsew signal input
flabel metal3 s 40300 616076 40600 616142 0 FreeSans 320 0 0 0 gpio6_1_in
port 1981 nsew signal output
flabel metal3 s 40300 615927 40600 615993 0 FreeSans 320 0 0 0 gpio6_1_hld_h_n
port 1982 nsew signal input
flabel metal3 s 40300 613754 40600 613820 0 FreeSans 320 0 0 0 gpio6_1_enable_vdda_h
port 1983 nsew signal input
flabel metal3 s 40300 613623 40600 613689 0 FreeSans 320 0 0 0 gpio6_1_analog_en
port 1984 nsew signal input
flabel metal3 s 40300 613422 40600 613488 0 FreeSans 320 0 0 0 gpio6_1_enable_inp_h
port 1985 nsew signal input
flabel metal3 s 40300 613153 40600 613273 0 FreeSans 320 0 0 0 gpio6_1_enable_vswitch_h
port 1986 nsew signal input
flabel metal3 s 40300 612577 40600 612697 0 FreeSans 320 0 0 0 gpio6_1_pad_a_noesd_h
port 1987 nsew signal bidirectional
flabel metal3 s 40300 612321 40600 612440 0 FreeSans 320 0 0 0 gpio6_1_pad_a_esd_0_h
port 1988 nsew signal bidirectional
flabel metal3 s 40300 612066 40600 612186 0 FreeSans 320 0 0 0 gpio6_1_pad_a_esd_1_h
port 1989 nsew signal bidirectional
flabel metal3 s 40300 641802 40600 641872 0 FreeSans 320 0 0 0 gpio6_1_zero
port 1990 nsew signal output
flabel metal3 s 40300 642252 40600 642322 0 FreeSans 320 0 0 0 gpio6_1_one
port 1991 nsew signal output
flabel metal3 s 40300 604995 40600 605061 0 FreeSans 320 0 0 0 gpio6_2_tie_hi_esd
port 1992 nsew signal output
flabel metal3 s 40300 600679 40600 600745 0 FreeSans 320 0 0 0 gpio6_2_dm[2]
port 1993 nsew signal input
flabel metal3 s 40300 604655 40600 604721 0 FreeSans 320 0 0 0 gpio6_2_dm[1]
port 1994 nsew signal input
flabel metal3 s 40300 604825 40600 604891 0 FreeSans 320 0 0 0 gpio6_2_dm[0]
port 1995 nsew signal input
flabel metal3 s 40300 604028 40600 604094 0 FreeSans 320 0 0 0 gpio6_2_slow
port 1996 nsew signal input
flabel metal3 s 40300 603889 40600 603955 0 FreeSans 320 0 0 0 gpio6_2_oe_n
port 1997 nsew signal input
flabel metal3 s 40300 602058 40600 602178 0 FreeSans 320 0 0 0 gpio6_2_tie_lo_esd
port 1998 nsew signal output
flabel metal3 s 40300 600509 40600 600575 0 FreeSans 320 0 0 0 gpio6_2_inp_dis
port 1999 nsew signal input
flabel metal3 s 40300 598169 40600 598243 0 FreeSans 320 0 0 0 gpio6_2_enable_vddio
port 2000 nsew signal input
flabel metal3 s 40300 596533 40600 596599 0 FreeSans 320 0 0 0 gpio6_2_vtrip_sel
port 2001 nsew signal input
flabel metal3 s 40300 592387 40600 592453 0 FreeSans 320 0 0 0 gpio6_2_ib_mode_sel[1]
port 2002 nsew signal input
flabel metal3 s 40300 596363 40600 596429 0 FreeSans 320 0 0 0 gpio6_2_ib_mode_sel[0]
port 2003 nsew signal input
flabel metal3 s 40300 593825 40600 593891 0 FreeSans 320 0 0 0 gpio6_2_out
port 2004 nsew signal input
flabel metal3 s 40300 588241 40600 588307 0 FreeSans 320 0 0 0 gpio6_2_slew_ctl[1]
port 2005 nsew signal input
flabel metal3 s 40300 592217 40600 592283 0 FreeSans 320 0 0 0 gpio6_2_slew_ctl[0]
port 2006 nsew signal input
flabel metal3 s 40300 592047 40600 592113 0 FreeSans 320 0 0 0 gpio6_2_analog_pol
port 2007 nsew signal input
flabel metal3 s 40300 589331 40600 589397 0 FreeSans 320 0 0 0 gpio6_2_analog_sel
port 2008 nsew signal input
flabel metal3 s 40300 588071 40600 588137 0 FreeSans 320 0 0 0 gpio6_2_hys_trim
port 2009 nsew signal input
flabel metal3 s 40300 587807 40600 587873 0 FreeSans 320 0 0 0 gpio6_2_vinref
port 2010 nsew signal input
flabel metal3 s 40300 584471 40600 584537 0 FreeSans 320 0 0 0 gpio6_2_hld_ovr
port 2011 nsew signal input
flabel metal3 s 40300 583876 40600 583942 0 FreeSans 320 0 0 0 gpio6_2_in_h
port 2012 nsew signal output
flabel metal3 s 40300 583427 40600 583493 0 FreeSans 320 0 0 0 gpio6_2_enable_h
port 2013 nsew signal input
flabel metal3 s 40300 583076 40600 583142 0 FreeSans 320 0 0 0 gpio6_2_in
port 2014 nsew signal output
flabel metal3 s 40300 582927 40600 582993 0 FreeSans 320 0 0 0 gpio6_2_hld_h_n
port 2015 nsew signal input
flabel metal3 s 40300 580754 40600 580820 0 FreeSans 320 0 0 0 gpio6_2_enable_vdda_h
port 2016 nsew signal input
flabel metal3 s 40300 580623 40600 580689 0 FreeSans 320 0 0 0 gpio6_2_analog_en
port 2017 nsew signal input
flabel metal3 s 40300 580422 40600 580488 0 FreeSans 320 0 0 0 gpio6_2_enable_inp_h
port 2018 nsew signal input
flabel metal3 s 40300 580153 40600 580273 0 FreeSans 320 0 0 0 gpio6_2_enable_vswitch_h
port 2019 nsew signal input
flabel metal3 s 40300 579577 40600 579697 0 FreeSans 320 0 0 0 gpio6_2_pad_a_noesd_h
port 2020 nsew signal bidirectional
flabel metal3 s 40300 579321 40600 579440 0 FreeSans 320 0 0 0 gpio6_2_pad_a_esd_0_h
port 2021 nsew signal bidirectional
flabel metal3 s 40300 579066 40600 579186 0 FreeSans 320 0 0 0 gpio6_2_pad_a_esd_1_h
port 2022 nsew signal bidirectional
flabel metal3 s 40300 608802 40600 608872 0 FreeSans 320 0 0 0 gpio6_2_zero
port 2023 nsew signal output
flabel metal3 s 40300 609252 40600 609322 0 FreeSans 320 0 0 0 gpio6_2_one
port 2024 nsew signal output
flabel metal3 s 40300 571995 40600 572061 0 FreeSans 320 0 0 0 gpio6_3_tie_hi_esd
port 2025 nsew signal output
flabel metal3 s 40300 567679 40600 567745 0 FreeSans 320 0 0 0 gpio6_3_dm[2]
port 2026 nsew signal input
flabel metal3 s 40300 571655 40600 571721 0 FreeSans 320 0 0 0 gpio6_3_dm[1]
port 2027 nsew signal input
flabel metal3 s 40300 571825 40600 571891 0 FreeSans 320 0 0 0 gpio6_3_dm[0]
port 2028 nsew signal input
flabel metal3 s 40300 571028 40600 571094 0 FreeSans 320 0 0 0 gpio6_3_slow
port 2029 nsew signal input
flabel metal3 s 40300 570889 40600 570955 0 FreeSans 320 0 0 0 gpio6_3_oe_n
port 2030 nsew signal input
flabel metal3 s 40300 569058 40600 569178 0 FreeSans 320 0 0 0 gpio6_3_tie_lo_esd
port 2031 nsew signal output
flabel metal3 s 40300 567509 40600 567575 0 FreeSans 320 0 0 0 gpio6_3_inp_dis
port 2032 nsew signal input
flabel metal3 s 40300 565169 40600 565243 0 FreeSans 320 0 0 0 gpio6_3_enable_vddio
port 2033 nsew signal input
flabel metal3 s 40300 563533 40600 563599 0 FreeSans 320 0 0 0 gpio6_3_vtrip_sel
port 2034 nsew signal input
flabel metal3 s 40300 559387 40600 559453 0 FreeSans 320 0 0 0 gpio6_3_ib_mode_sel[1]
port 2035 nsew signal input
flabel metal3 s 40300 563363 40600 563429 0 FreeSans 320 0 0 0 gpio6_3_ib_mode_sel[0]
port 2036 nsew signal input
flabel metal3 s 40300 560825 40600 560891 0 FreeSans 320 0 0 0 gpio6_3_out
port 2037 nsew signal input
flabel metal3 s 40300 555241 40600 555307 0 FreeSans 320 0 0 0 gpio6_3_slew_ctl[1]
port 2038 nsew signal input
flabel metal3 s 40300 559217 40600 559283 0 FreeSans 320 0 0 0 gpio6_3_slew_ctl[0]
port 2039 nsew signal input
flabel metal3 s 40300 559047 40600 559113 0 FreeSans 320 0 0 0 gpio6_3_analog_pol
port 2040 nsew signal input
flabel metal3 s 40300 556331 40600 556397 0 FreeSans 320 0 0 0 gpio6_3_analog_sel
port 2041 nsew signal input
flabel metal3 s 40300 555071 40600 555137 0 FreeSans 320 0 0 0 gpio6_3_hys_trim
port 2042 nsew signal input
flabel metal3 s 40300 554807 40600 554873 0 FreeSans 320 0 0 0 gpio6_3_vinref
port 2043 nsew signal input
flabel metal3 s 40300 551471 40600 551537 0 FreeSans 320 0 0 0 gpio6_3_hld_ovr
port 2044 nsew signal input
flabel metal3 s 40300 550876 40600 550942 0 FreeSans 320 0 0 0 gpio6_3_in_h
port 2045 nsew signal output
flabel metal3 s 40300 550427 40600 550493 0 FreeSans 320 0 0 0 gpio6_3_enable_h
port 2046 nsew signal input
flabel metal3 s 40300 550076 40600 550142 0 FreeSans 320 0 0 0 gpio6_3_in
port 2047 nsew signal output
flabel metal3 s 40300 549927 40600 549993 0 FreeSans 320 0 0 0 gpio6_3_hld_h_n
port 2048 nsew signal input
flabel metal3 s 40300 547754 40600 547820 0 FreeSans 320 0 0 0 gpio6_3_enable_vdda_h
port 2049 nsew signal input
flabel metal3 s 40300 547623 40600 547689 0 FreeSans 320 0 0 0 gpio6_3_analog_en
port 2050 nsew signal input
flabel metal3 s 40300 547422 40600 547488 0 FreeSans 320 0 0 0 gpio6_3_enable_inp_h
port 2051 nsew signal input
flabel metal3 s 40300 547153 40600 547273 0 FreeSans 320 0 0 0 gpio6_3_enable_vswitch_h
port 2052 nsew signal input
flabel metal3 s 40300 546577 40600 546697 0 FreeSans 320 0 0 0 gpio6_3_pad_a_noesd_h
port 2053 nsew signal bidirectional
flabel metal3 s 40300 546321 40600 546440 0 FreeSans 320 0 0 0 gpio6_3_pad_a_esd_0_h
port 2054 nsew signal bidirectional
flabel metal3 s 40300 546066 40600 546186 0 FreeSans 320 0 0 0 gpio6_3_pad_a_esd_1_h
port 2055 nsew signal bidirectional
flabel metal3 s 40300 575802 40600 575872 0 FreeSans 320 0 0 0 gpio6_3_zero
port 2056 nsew signal output
flabel metal3 s 40300 576252 40600 576322 0 FreeSans 320 0 0 0 gpio6_3_one
port 2057 nsew signal output
flabel metal3 s 40300 518895 40600 519295 0 FreeSans 320 0 0 0 vcap_w_cpos
port 2058 nsew signal bidirectional
flabel metal3 s 40600 514476 40900 514536 0 FreeSans 320 0 0 0 vref_w_ref_sel[1]
port 2059 nsew signal input
flabel metal3 s 40600 513495 40900 513555 0 FreeSans 320 0 0 0 vref_w_ref_sel[0]
port 2060 nsew signal input
flabel metal3 s 40600 508897 40900 509025 0 FreeSans 320 0 0 0 vref_w_vinref
port 2061 nsew signal output
flabel metal3 s 40600 508141 40900 508201 0 FreeSans 320 0 0 0 vref_w_ref_sel[2]
port 2062 nsew signal input
flabel metal3 s 40600 507943 40900 508003 0 FreeSans 320 0 0 0 vref_w_enable_h
port 2063 nsew signal input
flabel metal3 s 40600 507743 40900 507803 0 FreeSans 320 0 0 0 vref_w_hld_h_n
port 2064 nsew signal input
flabel metal3 s 40600 507455 40900 507515 0 FreeSans 320 0 0 0 vref_w_vrefgen_en
port 2065 nsew signal input
flabel metal3 s 40600 502627 40900 502687 0 FreeSans 320 0 0 0 vref_w_ref_sel[4]
port 2066 nsew signal input
flabel metal3 s 40600 502375 40900 502435 0 FreeSans 320 0 0 0 vref_w_ref_sel[3]
port 2067 nsew signal input
flabel metal3 s 40300 474395 40600 474461 0 FreeSans 320 0 0 0 gpio6_4_tie_hi_esd
port 2068 nsew signal output
flabel metal3 s 40300 470079 40600 470145 0 FreeSans 320 0 0 0 gpio6_4_dm[2]
port 2069 nsew signal input
flabel metal3 s 40300 474055 40600 474121 0 FreeSans 320 0 0 0 gpio6_4_dm[1]
port 2070 nsew signal input
flabel metal3 s 40300 474225 40600 474291 0 FreeSans 320 0 0 0 gpio6_4_dm[0]
port 2071 nsew signal input
flabel metal3 s 40300 473428 40600 473494 0 FreeSans 320 0 0 0 gpio6_4_slow
port 2072 nsew signal input
flabel metal3 s 40300 473289 40600 473355 0 FreeSans 320 0 0 0 gpio6_4_oe_n
port 2073 nsew signal input
flabel metal3 s 40300 471458 40600 471578 0 FreeSans 320 0 0 0 gpio6_4_tie_lo_esd
port 2074 nsew signal output
flabel metal3 s 40300 469909 40600 469975 0 FreeSans 320 0 0 0 gpio6_4_inp_dis
port 2075 nsew signal input
flabel metal3 s 40300 467569 40600 467643 0 FreeSans 320 0 0 0 gpio6_4_enable_vddio
port 2076 nsew signal input
flabel metal3 s 40300 465933 40600 465999 0 FreeSans 320 0 0 0 gpio6_4_vtrip_sel
port 2077 nsew signal input
flabel metal3 s 40300 461787 40600 461853 0 FreeSans 320 0 0 0 gpio6_4_ib_mode_sel[1]
port 2078 nsew signal input
flabel metal3 s 40300 465763 40600 465829 0 FreeSans 320 0 0 0 gpio6_4_ib_mode_sel[0]
port 2079 nsew signal input
flabel metal3 s 40300 463225 40600 463291 0 FreeSans 320 0 0 0 gpio6_4_out
port 2080 nsew signal input
flabel metal3 s 40300 457641 40600 457707 0 FreeSans 320 0 0 0 gpio6_4_slew_ctl[1]
port 2081 nsew signal input
flabel metal3 s 40300 461617 40600 461683 0 FreeSans 320 0 0 0 gpio6_4_slew_ctl[0]
port 2082 nsew signal input
flabel metal3 s 40300 461447 40600 461513 0 FreeSans 320 0 0 0 gpio6_4_analog_pol
port 2083 nsew signal input
flabel metal3 s 40300 458731 40600 458797 0 FreeSans 320 0 0 0 gpio6_4_analog_sel
port 2084 nsew signal input
flabel metal3 s 40300 457471 40600 457537 0 FreeSans 320 0 0 0 gpio6_4_hys_trim
port 2085 nsew signal input
flabel metal3 s 40300 457207 40600 457273 0 FreeSans 320 0 0 0 gpio6_4_vinref
port 2086 nsew signal input
flabel metal3 s 40300 453871 40600 453937 0 FreeSans 320 0 0 0 gpio6_4_hld_ovr
port 2087 nsew signal input
flabel metal3 s 40300 453276 40600 453342 0 FreeSans 320 0 0 0 gpio6_4_in_h
port 2088 nsew signal output
flabel metal3 s 40300 452827 40600 452893 0 FreeSans 320 0 0 0 gpio6_4_enable_h
port 2089 nsew signal input
flabel metal3 s 40300 452476 40600 452542 0 FreeSans 320 0 0 0 gpio6_4_in
port 2090 nsew signal output
flabel metal3 s 40300 452327 40600 452393 0 FreeSans 320 0 0 0 gpio6_4_hld_h_n
port 2091 nsew signal input
flabel metal3 s 40300 450154 40600 450220 0 FreeSans 320 0 0 0 gpio6_4_enable_vdda_h
port 2092 nsew signal input
flabel metal3 s 40300 450023 40600 450089 0 FreeSans 320 0 0 0 gpio6_4_analog_en
port 2093 nsew signal input
flabel metal3 s 40300 449822 40600 449888 0 FreeSans 320 0 0 0 gpio6_4_enable_inp_h
port 2094 nsew signal input
flabel metal3 s 40300 449553 40600 449673 0 FreeSans 320 0 0 0 gpio6_4_enable_vswitch_h
port 2095 nsew signal input
flabel metal3 s 40300 448977 40600 449097 0 FreeSans 320 0 0 0 gpio6_4_pad_a_noesd_h
port 2096 nsew signal bidirectional
flabel metal3 s 40300 448721 40600 448840 0 FreeSans 320 0 0 0 gpio6_4_pad_a_esd_0_h
port 2097 nsew signal bidirectional
flabel metal3 s 40300 448466 40600 448586 0 FreeSans 320 0 0 0 gpio6_4_pad_a_esd_1_h
port 2098 nsew signal bidirectional
flabel metal3 s 40300 478202 40600 478272 0 FreeSans 320 0 0 0 gpio6_4_zero
port 2099 nsew signal output
flabel metal3 s 40300 478652 40600 478722 0 FreeSans 320 0 0 0 gpio6_4_one
port 2100 nsew signal output
flabel metal3 s 40300 441395 40600 441461 0 FreeSans 320 0 0 0 gpio6_5_tie_hi_esd
port 2101 nsew signal output
flabel metal3 s 40300 437079 40600 437145 0 FreeSans 320 0 0 0 gpio6_5_dm[2]
port 2102 nsew signal input
flabel metal3 s 40300 441055 40600 441121 0 FreeSans 320 0 0 0 gpio6_5_dm[1]
port 2103 nsew signal input
flabel metal3 s 40300 441225 40600 441291 0 FreeSans 320 0 0 0 gpio6_5_dm[0]
port 2104 nsew signal input
flabel metal3 s 40300 440428 40600 440494 0 FreeSans 320 0 0 0 gpio6_5_slow
port 2105 nsew signal input
flabel metal3 s 40300 440289 40600 440355 0 FreeSans 320 0 0 0 gpio6_5_oe_n
port 2106 nsew signal input
flabel metal3 s 40300 438458 40600 438578 0 FreeSans 320 0 0 0 gpio6_5_tie_lo_esd
port 2107 nsew signal output
flabel metal3 s 40300 436909 40600 436975 0 FreeSans 320 0 0 0 gpio6_5_inp_dis
port 2108 nsew signal input
flabel metal3 s 40300 434569 40600 434643 0 FreeSans 320 0 0 0 gpio6_5_enable_vddio
port 2109 nsew signal input
flabel metal3 s 40300 432933 40600 432999 0 FreeSans 320 0 0 0 gpio6_5_vtrip_sel
port 2110 nsew signal input
flabel metal3 s 40300 428787 40600 428853 0 FreeSans 320 0 0 0 gpio6_5_ib_mode_sel[1]
port 2111 nsew signal input
flabel metal3 s 40300 432763 40600 432829 0 FreeSans 320 0 0 0 gpio6_5_ib_mode_sel[0]
port 2112 nsew signal input
flabel metal3 s 40300 430225 40600 430291 0 FreeSans 320 0 0 0 gpio6_5_out
port 2113 nsew signal input
flabel metal3 s 40300 424641 40600 424707 0 FreeSans 320 0 0 0 gpio6_5_slew_ctl[1]
port 2114 nsew signal input
flabel metal3 s 40300 428617 40600 428683 0 FreeSans 320 0 0 0 gpio6_5_slew_ctl[0]
port 2115 nsew signal input
flabel metal3 s 40300 428447 40600 428513 0 FreeSans 320 0 0 0 gpio6_5_analog_pol
port 2116 nsew signal input
flabel metal3 s 40300 425731 40600 425797 0 FreeSans 320 0 0 0 gpio6_5_analog_sel
port 2117 nsew signal input
flabel metal3 s 40300 424471 40600 424537 0 FreeSans 320 0 0 0 gpio6_5_hys_trim
port 2118 nsew signal input
flabel metal3 s 40300 424207 40600 424273 0 FreeSans 320 0 0 0 gpio6_5_vinref
port 2119 nsew signal input
flabel metal3 s 40300 420871 40600 420937 0 FreeSans 320 0 0 0 gpio6_5_hld_ovr
port 2120 nsew signal input
flabel metal3 s 40300 420276 40600 420342 0 FreeSans 320 0 0 0 gpio6_5_in_h
port 2121 nsew signal output
flabel metal3 s 40300 419827 40600 419893 0 FreeSans 320 0 0 0 gpio6_5_enable_h
port 2122 nsew signal input
flabel metal3 s 40300 419476 40600 419542 0 FreeSans 320 0 0 0 gpio6_5_in
port 2123 nsew signal output
flabel metal3 s 40300 419327 40600 419393 0 FreeSans 320 0 0 0 gpio6_5_hld_h_n
port 2124 nsew signal input
flabel metal3 s 40300 417154 40600 417220 0 FreeSans 320 0 0 0 gpio6_5_enable_vdda_h
port 2125 nsew signal input
flabel metal3 s 40300 417023 40600 417089 0 FreeSans 320 0 0 0 gpio6_5_analog_en
port 2126 nsew signal input
flabel metal3 s 40300 416822 40600 416888 0 FreeSans 320 0 0 0 gpio6_5_enable_inp_h
port 2127 nsew signal input
flabel metal3 s 40300 416553 40600 416673 0 FreeSans 320 0 0 0 gpio6_5_enable_vswitch_h
port 2128 nsew signal input
flabel metal3 s 40300 415977 40600 416097 0 FreeSans 320 0 0 0 gpio6_5_pad_a_noesd_h
port 2129 nsew signal bidirectional
flabel metal3 s 40300 415721 40600 415840 0 FreeSans 320 0 0 0 gpio6_5_pad_a_esd_0_h
port 2130 nsew signal bidirectional
flabel metal3 s 40300 415466 40600 415586 0 FreeSans 320 0 0 0 gpio6_5_pad_a_esd_1_h
port 2131 nsew signal bidirectional
flabel metal3 s 40300 445202 40600 445272 0 FreeSans 320 0 0 0 gpio6_5_zero
port 2132 nsew signal output
flabel metal3 s 40300 445652 40600 445722 0 FreeSans 320 0 0 0 gpio6_5_one
port 2133 nsew signal output
flabel metal3 s 40300 408395 40600 408461 0 FreeSans 320 0 0 0 gpio6_6_tie_hi_esd
port 2134 nsew signal output
flabel metal3 s 40300 404079 40600 404145 0 FreeSans 320 0 0 0 gpio6_6_dm[2]
port 2135 nsew signal input
flabel metal3 s 40300 408055 40600 408121 0 FreeSans 320 0 0 0 gpio6_6_dm[1]
port 2136 nsew signal input
flabel metal3 s 40300 408225 40600 408291 0 FreeSans 320 0 0 0 gpio6_6_dm[0]
port 2137 nsew signal input
flabel metal3 s 40300 407428 40600 407494 0 FreeSans 320 0 0 0 gpio6_6_slow
port 2138 nsew signal input
flabel metal3 s 40300 407289 40600 407355 0 FreeSans 320 0 0 0 gpio6_6_oe_n
port 2139 nsew signal input
flabel metal3 s 40300 405458 40600 405578 0 FreeSans 320 0 0 0 gpio6_6_tie_lo_esd
port 2140 nsew signal output
flabel metal3 s 40300 403909 40600 403975 0 FreeSans 320 0 0 0 gpio6_6_inp_dis
port 2141 nsew signal input
flabel metal3 s 40300 401569 40600 401643 0 FreeSans 320 0 0 0 gpio6_6_enable_vddio
port 2142 nsew signal input
flabel metal3 s 40300 399933 40600 399999 0 FreeSans 320 0 0 0 gpio6_6_vtrip_sel
port 2143 nsew signal input
flabel metal3 s 40300 395787 40600 395853 0 FreeSans 320 0 0 0 gpio6_6_ib_mode_sel[1]
port 2144 nsew signal input
flabel metal3 s 40300 399763 40600 399829 0 FreeSans 320 0 0 0 gpio6_6_ib_mode_sel[0]
port 2145 nsew signal input
flabel metal3 s 40300 397225 40600 397291 0 FreeSans 320 0 0 0 gpio6_6_out
port 2146 nsew signal input
flabel metal3 s 40300 391641 40600 391707 0 FreeSans 320 0 0 0 gpio6_6_slew_ctl[1]
port 2147 nsew signal input
flabel metal3 s 40300 395617 40600 395683 0 FreeSans 320 0 0 0 gpio6_6_slew_ctl[0]
port 2148 nsew signal input
flabel metal3 s 40300 395447 40600 395513 0 FreeSans 320 0 0 0 gpio6_6_analog_pol
port 2149 nsew signal input
flabel metal3 s 40300 392731 40600 392797 0 FreeSans 320 0 0 0 gpio6_6_analog_sel
port 2150 nsew signal input
flabel metal3 s 40300 391471 40600 391537 0 FreeSans 320 0 0 0 gpio6_6_hys_trim
port 2151 nsew signal input
flabel metal3 s 40300 391207 40600 391273 0 FreeSans 320 0 0 0 gpio6_6_vinref
port 2152 nsew signal input
flabel metal3 s 40300 387871 40600 387937 0 FreeSans 320 0 0 0 gpio6_6_hld_ovr
port 2153 nsew signal input
flabel metal3 s 40300 387276 40600 387342 0 FreeSans 320 0 0 0 gpio6_6_in_h
port 2154 nsew signal output
flabel metal3 s 40300 386827 40600 386893 0 FreeSans 320 0 0 0 gpio6_6_enable_h
port 2155 nsew signal input
flabel metal3 s 40300 386476 40600 386542 0 FreeSans 320 0 0 0 gpio6_6_in
port 2156 nsew signal output
flabel metal3 s 40300 386327 40600 386393 0 FreeSans 320 0 0 0 gpio6_6_hld_h_n
port 2157 nsew signal input
flabel metal3 s 40300 384154 40600 384220 0 FreeSans 320 0 0 0 gpio6_6_enable_vdda_h
port 2158 nsew signal input
flabel metal3 s 40300 384023 40600 384089 0 FreeSans 320 0 0 0 gpio6_6_analog_en
port 2159 nsew signal input
flabel metal3 s 40300 383822 40600 383888 0 FreeSans 320 0 0 0 gpio6_6_enable_inp_h
port 2160 nsew signal input
flabel metal3 s 40300 383553 40600 383673 0 FreeSans 320 0 0 0 gpio6_6_enable_vswitch_h
port 2161 nsew signal input
flabel metal3 s 40300 382977 40600 383097 0 FreeSans 320 0 0 0 gpio6_6_pad_a_noesd_h
port 2162 nsew signal bidirectional
flabel metal3 s 40300 382721 40600 382840 0 FreeSans 320 0 0 0 gpio6_6_pad_a_esd_0_h
port 2163 nsew signal bidirectional
flabel metal3 s 40300 382466 40600 382586 0 FreeSans 320 0 0 0 gpio6_6_pad_a_esd_1_h
port 2164 nsew signal bidirectional
flabel metal3 s 40300 412202 40600 412272 0 FreeSans 320 0 0 0 gpio6_6_zero
port 2165 nsew signal output
flabel metal3 s 40300 412652 40600 412722 0 FreeSans 320 0 0 0 gpio6_6_one
port 2166 nsew signal output
flabel metal3 s 40300 375395 40600 375461 0 FreeSans 320 0 0 0 gpio6_7_tie_hi_esd
port 2167 nsew signal output
flabel metal3 s 40300 371079 40600 371145 0 FreeSans 320 0 0 0 gpio6_7_dm[2]
port 2168 nsew signal input
flabel metal3 s 40300 375055 40600 375121 0 FreeSans 320 0 0 0 gpio6_7_dm[1]
port 2169 nsew signal input
flabel metal3 s 40300 375225 40600 375291 0 FreeSans 320 0 0 0 gpio6_7_dm[0]
port 2170 nsew signal input
flabel metal3 s 40300 374428 40600 374494 0 FreeSans 320 0 0 0 gpio6_7_slow
port 2171 nsew signal input
flabel metal3 s 40300 374289 40600 374355 0 FreeSans 320 0 0 0 gpio6_7_oe_n
port 2172 nsew signal input
flabel metal3 s 40300 372458 40600 372578 0 FreeSans 320 0 0 0 gpio6_7_tie_lo_esd
port 2173 nsew signal output
flabel metal3 s 40300 370909 40600 370975 0 FreeSans 320 0 0 0 gpio6_7_inp_dis
port 2174 nsew signal input
flabel metal3 s 40300 368569 40600 368643 0 FreeSans 320 0 0 0 gpio6_7_enable_vddio
port 2175 nsew signal input
flabel metal3 s 40300 366933 40600 366999 0 FreeSans 320 0 0 0 gpio6_7_vtrip_sel
port 2176 nsew signal input
flabel metal3 s 40300 362787 40600 362853 0 FreeSans 320 0 0 0 gpio6_7_ib_mode_sel[1]
port 2177 nsew signal input
flabel metal3 s 40300 366763 40600 366829 0 FreeSans 320 0 0 0 gpio6_7_ib_mode_sel[0]
port 2178 nsew signal input
flabel metal3 s 40300 364225 40600 364291 0 FreeSans 320 0 0 0 gpio6_7_out
port 2179 nsew signal input
flabel metal3 s 40300 358641 40600 358707 0 FreeSans 320 0 0 0 gpio6_7_slew_ctl[1]
port 2180 nsew signal input
flabel metal3 s 40300 362617 40600 362683 0 FreeSans 320 0 0 0 gpio6_7_slew_ctl[0]
port 2181 nsew signal input
flabel metal3 s 40300 362447 40600 362513 0 FreeSans 320 0 0 0 gpio6_7_analog_pol
port 2182 nsew signal input
flabel metal3 s 40300 359731 40600 359797 0 FreeSans 320 0 0 0 gpio6_7_analog_sel
port 2183 nsew signal input
flabel metal3 s 40300 358471 40600 358537 0 FreeSans 320 0 0 0 gpio6_7_hys_trim
port 2184 nsew signal input
flabel metal3 s 40300 358207 40600 358273 0 FreeSans 320 0 0 0 gpio6_7_vinref
port 2185 nsew signal input
flabel metal3 s 40300 354871 40600 354937 0 FreeSans 320 0 0 0 gpio6_7_hld_ovr
port 2186 nsew signal input
flabel metal3 s 40300 354276 40600 354342 0 FreeSans 320 0 0 0 gpio6_7_in_h
port 2187 nsew signal output
flabel metal3 s 40300 353827 40600 353893 0 FreeSans 320 0 0 0 gpio6_7_enable_h
port 2188 nsew signal input
flabel metal3 s 40300 353476 40600 353542 0 FreeSans 320 0 0 0 gpio6_7_in
port 2189 nsew signal output
flabel metal3 s 40300 353327 40600 353393 0 FreeSans 320 0 0 0 gpio6_7_hld_h_n
port 2190 nsew signal input
flabel metal3 s 40300 351154 40600 351220 0 FreeSans 320 0 0 0 gpio6_7_enable_vdda_h
port 2191 nsew signal input
flabel metal3 s 40300 351023 40600 351089 0 FreeSans 320 0 0 0 gpio6_7_analog_en
port 2192 nsew signal input
flabel metal3 s 40300 350822 40600 350888 0 FreeSans 320 0 0 0 gpio6_7_enable_inp_h
port 2193 nsew signal input
flabel metal3 s 40300 350553 40600 350673 0 FreeSans 320 0 0 0 gpio6_7_enable_vswitch_h
port 2194 nsew signal input
flabel metal3 s 40300 349977 40600 350097 0 FreeSans 320 0 0 0 gpio6_7_pad_a_noesd_h
port 2195 nsew signal bidirectional
flabel metal3 s 40300 349721 40600 349840 0 FreeSans 320 0 0 0 gpio6_7_pad_a_esd_0_h
port 2196 nsew signal bidirectional
flabel metal3 s 40300 349466 40600 349586 0 FreeSans 320 0 0 0 gpio6_7_pad_a_esd_1_h
port 2197 nsew signal bidirectional
flabel metal3 s 40300 379202 40600 379272 0 FreeSans 320 0 0 0 gpio6_7_zero
port 2198 nsew signal output
flabel metal3 s 40300 379652 40600 379722 0 FreeSans 320 0 0 0 gpio6_7_one
port 2199 nsew signal output
flabel metal3 s 40542 282002 40842 282072 0 FreeSans 320 0 0 0 gpio7_0_tie_lo_esd
port 2200 nsew signal output
flabel metal3 s 40538 281424 40838 281494 0 FreeSans 320 0 0 0 gpio7_0_in
port 2201 nsew signal output
flabel metal3 s 40542 281704 40842 281774 0 FreeSans 320 0 0 0 gpio7_0_tie_hi_esd
port 2202 nsew signal output
flabel metal3 s 40542 281112 40842 281182 0 FreeSans 320 0 0 0 gpio7_0_enable_vddio
port 2203 nsew signal input
flabel metal3 s 40542 280838 40842 280908 0 FreeSans 320 0 0 0 gpio7_0_slow
port 2204 nsew signal input
flabel metal3 s 40542 280490 40842 280618 0 FreeSans 320 0 0 0 gpio7_0_pad_a_esd_0_h
port 2205 nsew signal bidirectional
flabel metal3 s 40542 279058 40842 279188 0 FreeSans 320 0 0 0 gpio7_0_pad_a_esd_1_h
port 2206 nsew signal bidirectional
flabel metal3 s 40542 277964 40842 278178 0 FreeSans 320 0 0 0 gpio7_0_pad_a_noesd_h
port 2207 nsew signal bidirectional
flabel metal3 s 40542 277332 40842 277402 0 FreeSans 320 0 0 0 gpio7_0_analog_en
port 2208 nsew signal input
flabel metal3 s 40542 274572 40842 274642 0 FreeSans 320 0 0 0 gpio7_0_analog_pol
port 2209 nsew signal input
flabel metal3 s 40542 273992 40842 274062 0 FreeSans 320 0 0 0 gpio7_0_inp_dis
port 2210 nsew signal input
flabel metal3 s 40542 272826 40842 272896 0 FreeSans 320 0 0 0 gpio7_0_enable_inp_h
port 2211 nsew signal input
flabel metal3 s 40542 272370 40842 272440 0 FreeSans 320 0 0 0 gpio7_0_enable_h
port 2212 nsew signal input
flabel metal3 s 40542 271916 40842 271986 0 FreeSans 320 0 0 0 gpio7_0_hld_h_n
port 2213 nsew signal input
flabel metal3 s 40542 271298 40842 271368 0 FreeSans 320 0 0 0 gpio7_0_analog_sel
port 2214 nsew signal input
flabel metal3 s 40542 270854 40842 270924 0 FreeSans 320 0 0 0 gpio7_0_dm[2]
port 2215 nsew signal input
flabel metal3 s 40542 278528 40842 278598 0 FreeSans 320 0 0 0 gpio7_0_dm[1]
port 2216 nsew signal input
flabel metal3 s 40542 275120 40842 275190 0 FreeSans 320 0 0 0 gpio7_0_dm[0]
port 2217 nsew signal input
flabel metal3 s 40542 270370 40842 270440 0 FreeSans 320 0 0 0 gpio7_0_hld_ovr
port 2218 nsew signal input
flabel metal3 s 40542 269598 40842 269668 0 FreeSans 320 0 0 0 gpio7_0_out
port 2219 nsew signal input
flabel metal3 s 40542 268398 40842 268468 0 FreeSans 320 0 0 0 gpio7_0_enable_vswitch_h
port 2220 nsew signal input
flabel metal3 s 40542 267678 40842 267748 0 FreeSans 320 0 0 0 gpio7_0_enable_vdda_h
port 2221 nsew signal input
flabel metal3 s 40542 266816 40842 266886 0 FreeSans 320 0 0 0 gpio7_0_vtrip_sel
port 2222 nsew signal input
flabel metal3 s 40542 266472 40842 266542 0 FreeSans 320 0 0 0 gpio7_0_ib_mode_sel
port 2223 nsew signal input
flabel metal3 s 40542 266062 40842 266132 0 FreeSans 320 0 0 0 gpio7_0_oe_n
port 2224 nsew signal input
flabel metal3 s 40542 265480 40842 265604 0 FreeSans 320 0 0 0 gpio7_0_in_h
port 2225 nsew signal output
flabel metal3 s 40542 283202 40842 283272 0 FreeSans 320 0 0 0 gpio7_0_zero
port 2226 nsew signal output
flabel metal3 s 40542 283652 40842 283722 0 FreeSans 320 0 0 0 gpio7_0_one
port 2227 nsew signal output
flabel metal3 s 40542 261002 40842 261072 0 FreeSans 320 0 0 0 gpio7_1_tie_lo_esd
port 2228 nsew signal output
flabel metal3 s 40538 260424 40838 260494 0 FreeSans 320 0 0 0 gpio7_1_in
port 2229 nsew signal output
flabel metal3 s 40542 260704 40842 260774 0 FreeSans 320 0 0 0 gpio7_1_tie_hi_esd
port 2230 nsew signal output
flabel metal3 s 40542 260112 40842 260182 0 FreeSans 320 0 0 0 gpio7_1_enable_vddio
port 2231 nsew signal input
flabel metal3 s 40542 259838 40842 259908 0 FreeSans 320 0 0 0 gpio7_1_slow
port 2232 nsew signal input
flabel metal3 s 40542 259490 40842 259618 0 FreeSans 320 0 0 0 gpio7_1_pad_a_esd_0_h
port 2233 nsew signal bidirectional
flabel metal3 s 40542 258058 40842 258188 0 FreeSans 320 0 0 0 gpio7_1_pad_a_esd_1_h
port 2234 nsew signal bidirectional
flabel metal3 s 40542 256964 40842 257178 0 FreeSans 320 0 0 0 gpio7_1_pad_a_noesd_h
port 2235 nsew signal bidirectional
flabel metal3 s 40542 256332 40842 256402 0 FreeSans 320 0 0 0 gpio7_1_analog_en
port 2236 nsew signal input
flabel metal3 s 40542 253572 40842 253642 0 FreeSans 320 0 0 0 gpio7_1_analog_pol
port 2237 nsew signal input
flabel metal3 s 40542 252992 40842 253062 0 FreeSans 320 0 0 0 gpio7_1_inp_dis
port 2238 nsew signal input
flabel metal3 s 40542 251826 40842 251896 0 FreeSans 320 0 0 0 gpio7_1_enable_inp_h
port 2239 nsew signal input
flabel metal3 s 40542 251370 40842 251440 0 FreeSans 320 0 0 0 gpio7_1_enable_h
port 2240 nsew signal input
flabel metal3 s 40542 250916 40842 250986 0 FreeSans 320 0 0 0 gpio7_1_hld_h_n
port 2241 nsew signal input
flabel metal3 s 40542 250298 40842 250368 0 FreeSans 320 0 0 0 gpio7_1_analog_sel
port 2242 nsew signal input
flabel metal3 s 40542 249854 40842 249924 0 FreeSans 320 0 0 0 gpio7_1_dm[2]
port 2243 nsew signal input
flabel metal3 s 40542 257528 40842 257598 0 FreeSans 320 0 0 0 gpio7_1_dm[1]
port 2244 nsew signal input
flabel metal3 s 40542 254120 40842 254190 0 FreeSans 320 0 0 0 gpio7_1_dm[0]
port 2245 nsew signal input
flabel metal3 s 40542 249370 40842 249440 0 FreeSans 320 0 0 0 gpio7_1_hld_ovr
port 2246 nsew signal input
flabel metal3 s 40542 248598 40842 248668 0 FreeSans 320 0 0 0 gpio7_1_out
port 2247 nsew signal input
flabel metal3 s 40542 247398 40842 247468 0 FreeSans 320 0 0 0 gpio7_1_enable_vswitch_h
port 2248 nsew signal input
flabel metal3 s 40542 246678 40842 246748 0 FreeSans 320 0 0 0 gpio7_1_enable_vdda_h
port 2249 nsew signal input
flabel metal3 s 40542 245816 40842 245886 0 FreeSans 320 0 0 0 gpio7_1_vtrip_sel
port 2250 nsew signal input
flabel metal3 s 40542 245472 40842 245542 0 FreeSans 320 0 0 0 gpio7_1_ib_mode_sel
port 2251 nsew signal input
flabel metal3 s 40542 245062 40842 245132 0 FreeSans 320 0 0 0 gpio7_1_oe_n
port 2252 nsew signal input
flabel metal3 s 40542 244480 40842 244604 0 FreeSans 320 0 0 0 gpio7_1_in_h
port 2253 nsew signal output
flabel metal3 s 40542 262202 40842 262272 0 FreeSans 320 0 0 0 gpio7_1_zero
port 2254 nsew signal output
flabel metal3 s 40542 262652 40842 262722 0 FreeSans 320 0 0 0 gpio7_1_one
port 2255 nsew signal output
flabel metal3 s 40542 240002 40842 240072 0 FreeSans 320 0 0 0 gpio7_2_tie_lo_esd
port 2256 nsew signal output
flabel metal3 s 40538 239424 40838 239494 0 FreeSans 320 0 0 0 gpio7_2_in
port 2257 nsew signal output
flabel metal3 s 40542 239704 40842 239774 0 FreeSans 320 0 0 0 gpio7_2_tie_hi_esd
port 2258 nsew signal output
flabel metal3 s 40542 239112 40842 239182 0 FreeSans 320 0 0 0 gpio7_2_enable_vddio
port 2259 nsew signal input
flabel metal3 s 40542 238838 40842 238908 0 FreeSans 320 0 0 0 gpio7_2_slow
port 2260 nsew signal input
flabel metal3 s 40542 238490 40842 238618 0 FreeSans 320 0 0 0 gpio7_2_pad_a_esd_0_h
port 2261 nsew signal bidirectional
flabel metal3 s 40542 237058 40842 237188 0 FreeSans 320 0 0 0 gpio7_2_pad_a_esd_1_h
port 2262 nsew signal bidirectional
flabel metal3 s 40542 235964 40842 236178 0 FreeSans 320 0 0 0 gpio7_2_pad_a_noesd_h
port 2263 nsew signal bidirectional
flabel metal3 s 40542 235332 40842 235402 0 FreeSans 320 0 0 0 gpio7_2_analog_en
port 2264 nsew signal input
flabel metal3 s 40542 232572 40842 232642 0 FreeSans 320 0 0 0 gpio7_2_analog_pol
port 2265 nsew signal input
flabel metal3 s 40542 231992 40842 232062 0 FreeSans 320 0 0 0 gpio7_2_inp_dis
port 2266 nsew signal input
flabel metal3 s 40542 230826 40842 230896 0 FreeSans 320 0 0 0 gpio7_2_enable_inp_h
port 2267 nsew signal input
flabel metal3 s 40542 230370 40842 230440 0 FreeSans 320 0 0 0 gpio7_2_enable_h
port 2268 nsew signal input
flabel metal3 s 40542 229916 40842 229986 0 FreeSans 320 0 0 0 gpio7_2_hld_h_n
port 2269 nsew signal input
flabel metal3 s 40542 229298 40842 229368 0 FreeSans 320 0 0 0 gpio7_2_analog_sel
port 2270 nsew signal input
flabel metal3 s 40542 228854 40842 228924 0 FreeSans 320 0 0 0 gpio7_2_dm[2]
port 2271 nsew signal input
flabel metal3 s 40542 236528 40842 236598 0 FreeSans 320 0 0 0 gpio7_2_dm[1]
port 2272 nsew signal input
flabel metal3 s 40542 233120 40842 233190 0 FreeSans 320 0 0 0 gpio7_2_dm[0]
port 2273 nsew signal input
flabel metal3 s 40542 228370 40842 228440 0 FreeSans 320 0 0 0 gpio7_2_hld_ovr
port 2274 nsew signal input
flabel metal3 s 40542 227598 40842 227668 0 FreeSans 320 0 0 0 gpio7_2_out
port 2275 nsew signal input
flabel metal3 s 40542 226398 40842 226468 0 FreeSans 320 0 0 0 gpio7_2_enable_vswitch_h
port 2276 nsew signal input
flabel metal3 s 40542 225678 40842 225748 0 FreeSans 320 0 0 0 gpio7_2_enable_vdda_h
port 2277 nsew signal input
flabel metal3 s 40542 224816 40842 224886 0 FreeSans 320 0 0 0 gpio7_2_vtrip_sel
port 2278 nsew signal input
flabel metal3 s 40542 224472 40842 224542 0 FreeSans 320 0 0 0 gpio7_2_ib_mode_sel
port 2279 nsew signal input
flabel metal3 s 40542 224062 40842 224132 0 FreeSans 320 0 0 0 gpio7_2_oe_n
port 2280 nsew signal input
flabel metal3 s 40542 223480 40842 223604 0 FreeSans 320 0 0 0 gpio7_2_in_h
port 2281 nsew signal output
flabel metal3 s 40542 241202 40842 241272 0 FreeSans 320 0 0 0 gpio7_2_zero
port 2282 nsew signal output
flabel metal3 s 40542 241652 40842 241722 0 FreeSans 320 0 0 0 gpio7_2_one
port 2283 nsew signal output
flabel metal3 s 40542 219002 40842 219072 0 FreeSans 320 0 0 0 gpio7_3_tie_lo_esd
port 2284 nsew signal output
flabel metal3 s 40538 218424 40838 218494 0 FreeSans 320 0 0 0 gpio7_3_in
port 2285 nsew signal output
flabel metal3 s 40542 218704 40842 218774 0 FreeSans 320 0 0 0 gpio7_3_tie_hi_esd
port 2286 nsew signal output
flabel metal3 s 40542 218112 40842 218182 0 FreeSans 320 0 0 0 gpio7_3_enable_vddio
port 2287 nsew signal input
flabel metal3 s 40542 217838 40842 217908 0 FreeSans 320 0 0 0 gpio7_3_slow
port 2288 nsew signal input
flabel metal3 s 40542 217490 40842 217618 0 FreeSans 320 0 0 0 gpio7_3_pad_a_esd_0_h
port 2289 nsew signal bidirectional
flabel metal3 s 40542 216058 40842 216188 0 FreeSans 320 0 0 0 gpio7_3_pad_a_esd_1_h
port 2290 nsew signal bidirectional
flabel metal3 s 40542 214964 40842 215178 0 FreeSans 320 0 0 0 gpio7_3_pad_a_noesd_h
port 2291 nsew signal bidirectional
flabel metal3 s 40542 214332 40842 214402 0 FreeSans 320 0 0 0 gpio7_3_analog_en
port 2292 nsew signal input
flabel metal3 s 40542 211572 40842 211642 0 FreeSans 320 0 0 0 gpio7_3_analog_pol
port 2293 nsew signal input
flabel metal3 s 40542 210992 40842 211062 0 FreeSans 320 0 0 0 gpio7_3_inp_dis
port 2294 nsew signal input
flabel metal3 s 40542 209826 40842 209896 0 FreeSans 320 0 0 0 gpio7_3_enable_inp_h
port 2295 nsew signal input
flabel metal3 s 40542 209370 40842 209440 0 FreeSans 320 0 0 0 gpio7_3_enable_h
port 2296 nsew signal input
flabel metal3 s 40542 208916 40842 208986 0 FreeSans 320 0 0 0 gpio7_3_hld_h_n
port 2297 nsew signal input
flabel metal3 s 40542 208298 40842 208368 0 FreeSans 320 0 0 0 gpio7_3_analog_sel
port 2298 nsew signal input
flabel metal3 s 40542 207854 40842 207924 0 FreeSans 320 0 0 0 gpio7_3_dm[2]
port 2299 nsew signal input
flabel metal3 s 40542 215528 40842 215598 0 FreeSans 320 0 0 0 gpio7_3_dm[1]
port 2300 nsew signal input
flabel metal3 s 40542 212120 40842 212190 0 FreeSans 320 0 0 0 gpio7_3_dm[0]
port 2301 nsew signal input
flabel metal3 s 40542 207370 40842 207440 0 FreeSans 320 0 0 0 gpio7_3_hld_ovr
port 2302 nsew signal input
flabel metal3 s 40542 206598 40842 206668 0 FreeSans 320 0 0 0 gpio7_3_out
port 2303 nsew signal input
flabel metal3 s 40542 205398 40842 205468 0 FreeSans 320 0 0 0 gpio7_3_enable_vswitch_h
port 2304 nsew signal input
flabel metal3 s 40542 204678 40842 204748 0 FreeSans 320 0 0 0 gpio7_3_enable_vdda_h
port 2305 nsew signal input
flabel metal3 s 40542 203816 40842 203886 0 FreeSans 320 0 0 0 gpio7_3_vtrip_sel
port 2306 nsew signal input
flabel metal3 s 40542 203472 40842 203542 0 FreeSans 320 0 0 0 gpio7_3_ib_mode_sel
port 2307 nsew signal input
flabel metal3 s 40542 203062 40842 203132 0 FreeSans 320 0 0 0 gpio7_3_oe_n
port 2308 nsew signal input
flabel metal3 s 40542 202480 40842 202604 0 FreeSans 320 0 0 0 gpio7_3_in_h
port 2309 nsew signal output
flabel metal3 s 40542 220202 40842 220272 0 FreeSans 320 0 0 0 gpio7_3_zero
port 2310 nsew signal output
flabel metal3 s 40542 220652 40842 220722 0 FreeSans 320 0 0 0 gpio7_3_one
port 2311 nsew signal output
flabel metal3 s 40542 155002 40842 155072 0 FreeSans 320 0 0 0 gpio7_4_tie_lo_esd
port 2312 nsew signal output
flabel metal3 s 40538 154424 40838 154494 0 FreeSans 320 0 0 0 gpio7_4_in
port 2313 nsew signal output
flabel metal3 s 40542 154704 40842 154774 0 FreeSans 320 0 0 0 gpio7_4_tie_hi_esd
port 2314 nsew signal output
flabel metal3 s 40542 154112 40842 154182 0 FreeSans 320 0 0 0 gpio7_4_enable_vddio
port 2315 nsew signal input
flabel metal3 s 40542 153838 40842 153908 0 FreeSans 320 0 0 0 gpio7_4_slow
port 2316 nsew signal input
flabel metal3 s 40542 153490 40842 153618 0 FreeSans 320 0 0 0 gpio7_4_pad_a_esd_0_h
port 2317 nsew signal bidirectional
flabel metal3 s 40542 152058 40842 152188 0 FreeSans 320 0 0 0 gpio7_4_pad_a_esd_1_h
port 2318 nsew signal bidirectional
flabel metal3 s 40542 150964 40842 151178 0 FreeSans 320 0 0 0 gpio7_4_pad_a_noesd_h
port 2319 nsew signal bidirectional
flabel metal3 s 40542 150332 40842 150402 0 FreeSans 320 0 0 0 gpio7_4_analog_en
port 2320 nsew signal input
flabel metal3 s 40542 147572 40842 147642 0 FreeSans 320 0 0 0 gpio7_4_analog_pol
port 2321 nsew signal input
flabel metal3 s 40542 146992 40842 147062 0 FreeSans 320 0 0 0 gpio7_4_inp_dis
port 2322 nsew signal input
flabel metal3 s 40542 145826 40842 145896 0 FreeSans 320 0 0 0 gpio7_4_enable_inp_h
port 2323 nsew signal input
flabel metal3 s 40542 145370 40842 145440 0 FreeSans 320 0 0 0 gpio7_4_enable_h
port 2324 nsew signal input
flabel metal3 s 40542 144916 40842 144986 0 FreeSans 320 0 0 0 gpio7_4_hld_h_n
port 2325 nsew signal input
flabel metal3 s 40542 144298 40842 144368 0 FreeSans 320 0 0 0 gpio7_4_analog_sel
port 2326 nsew signal input
flabel metal3 s 40542 143854 40842 143924 0 FreeSans 320 0 0 0 gpio7_4_dm[2]
port 2327 nsew signal input
flabel metal3 s 40542 151528 40842 151598 0 FreeSans 320 0 0 0 gpio7_4_dm[1]
port 2328 nsew signal input
flabel metal3 s 40542 148120 40842 148190 0 FreeSans 320 0 0 0 gpio7_4_dm[0]
port 2329 nsew signal input
flabel metal3 s 40542 143370 40842 143440 0 FreeSans 320 0 0 0 gpio7_4_hld_ovr
port 2330 nsew signal input
flabel metal3 s 40542 142598 40842 142668 0 FreeSans 320 0 0 0 gpio7_4_out
port 2331 nsew signal input
flabel metal3 s 40542 141398 40842 141468 0 FreeSans 320 0 0 0 gpio7_4_enable_vswitch_h
port 2332 nsew signal input
flabel metal3 s 40542 140678 40842 140748 0 FreeSans 320 0 0 0 gpio7_4_enable_vdda_h
port 2333 nsew signal input
flabel metal3 s 40542 139816 40842 139886 0 FreeSans 320 0 0 0 gpio7_4_vtrip_sel
port 2334 nsew signal input
flabel metal3 s 40542 139472 40842 139542 0 FreeSans 320 0 0 0 gpio7_4_ib_mode_sel
port 2335 nsew signal input
flabel metal3 s 40542 139062 40842 139132 0 FreeSans 320 0 0 0 gpio7_4_oe_n
port 2336 nsew signal input
flabel metal3 s 40542 138480 40842 138604 0 FreeSans 320 0 0 0 gpio7_4_in_h
port 2337 nsew signal output
flabel metal3 s 40542 156202 40842 156272 0 FreeSans 320 0 0 0 gpio7_4_zero
port 2338 nsew signal output
flabel metal3 s 40542 156652 40842 156722 0 FreeSans 320 0 0 0 gpio7_4_one
port 2339 nsew signal output
flabel metal3 s 40542 134002 40842 134072 0 FreeSans 320 0 0 0 gpio7_5_tie_lo_esd
port 2340 nsew signal output
flabel metal3 s 40538 133424 40838 133494 0 FreeSans 320 0 0 0 gpio7_5_in
port 2341 nsew signal output
flabel metal3 s 40542 133704 40842 133774 0 FreeSans 320 0 0 0 gpio7_5_tie_hi_esd
port 2342 nsew signal output
flabel metal3 s 40542 133112 40842 133182 0 FreeSans 320 0 0 0 gpio7_5_enable_vddio
port 2343 nsew signal input
flabel metal3 s 40542 132838 40842 132908 0 FreeSans 320 0 0 0 gpio7_5_slow
port 2344 nsew signal input
flabel metal3 s 40542 132490 40842 132618 0 FreeSans 320 0 0 0 gpio7_5_pad_a_esd_0_h
port 2345 nsew signal bidirectional
flabel metal3 s 40542 131058 40842 131188 0 FreeSans 320 0 0 0 gpio7_5_pad_a_esd_1_h
port 2346 nsew signal bidirectional
flabel metal3 s 40542 129964 40842 130178 0 FreeSans 320 0 0 0 gpio7_5_pad_a_noesd_h
port 2347 nsew signal bidirectional
flabel metal3 s 40542 129332 40842 129402 0 FreeSans 320 0 0 0 gpio7_5_analog_en
port 2348 nsew signal input
flabel metal3 s 40542 126572 40842 126642 0 FreeSans 320 0 0 0 gpio7_5_analog_pol
port 2349 nsew signal input
flabel metal3 s 40542 125992 40842 126062 0 FreeSans 320 0 0 0 gpio7_5_inp_dis
port 2350 nsew signal input
flabel metal3 s 40542 124826 40842 124896 0 FreeSans 320 0 0 0 gpio7_5_enable_inp_h
port 2351 nsew signal input
flabel metal3 s 40542 124370 40842 124440 0 FreeSans 320 0 0 0 gpio7_5_enable_h
port 2352 nsew signal input
flabel metal3 s 40542 123916 40842 123986 0 FreeSans 320 0 0 0 gpio7_5_hld_h_n
port 2353 nsew signal input
flabel metal3 s 40542 123298 40842 123368 0 FreeSans 320 0 0 0 gpio7_5_analog_sel
port 2354 nsew signal input
flabel metal3 s 40542 122854 40842 122924 0 FreeSans 320 0 0 0 gpio7_5_dm[2]
port 2355 nsew signal input
flabel metal3 s 40542 130528 40842 130598 0 FreeSans 320 0 0 0 gpio7_5_dm[1]
port 2356 nsew signal input
flabel metal3 s 40542 127120 40842 127190 0 FreeSans 320 0 0 0 gpio7_5_dm[0]
port 2357 nsew signal input
flabel metal3 s 40542 122370 40842 122440 0 FreeSans 320 0 0 0 gpio7_5_hld_ovr
port 2358 nsew signal input
flabel metal3 s 40542 121598 40842 121668 0 FreeSans 320 0 0 0 gpio7_5_out
port 2359 nsew signal input
flabel metal3 s 40542 120398 40842 120468 0 FreeSans 320 0 0 0 gpio7_5_enable_vswitch_h
port 2360 nsew signal input
flabel metal3 s 40542 119678 40842 119748 0 FreeSans 320 0 0 0 gpio7_5_enable_vdda_h
port 2361 nsew signal input
flabel metal3 s 40542 118816 40842 118886 0 FreeSans 320 0 0 0 gpio7_5_vtrip_sel
port 2362 nsew signal input
flabel metal3 s 40542 118472 40842 118542 0 FreeSans 320 0 0 0 gpio7_5_ib_mode_sel
port 2363 nsew signal input
flabel metal3 s 40542 118062 40842 118132 0 FreeSans 320 0 0 0 gpio7_5_oe_n
port 2364 nsew signal input
flabel metal3 s 40542 117480 40842 117604 0 FreeSans 320 0 0 0 gpio7_5_in_h
port 2365 nsew signal output
flabel metal3 s 40542 135202 40842 135272 0 FreeSans 320 0 0 0 gpio7_5_zero
port 2366 nsew signal output
flabel metal3 s 40542 135652 40842 135722 0 FreeSans 320 0 0 0 gpio7_5_one
port 2367 nsew signal output
flabel metal3 s 40542 113002 40842 113072 0 FreeSans 320 0 0 0 gpio7_6_tie_lo_esd
port 2368 nsew signal output
flabel metal3 s 40538 112424 40838 112494 0 FreeSans 320 0 0 0 gpio7_6_in
port 2369 nsew signal output
flabel metal3 s 40542 112704 40842 112774 0 FreeSans 320 0 0 0 gpio7_6_tie_hi_esd
port 2370 nsew signal output
flabel metal3 s 40542 112112 40842 112182 0 FreeSans 320 0 0 0 gpio7_6_enable_vddio
port 2371 nsew signal input
flabel metal3 s 40542 111838 40842 111908 0 FreeSans 320 0 0 0 gpio7_6_slow
port 2372 nsew signal input
flabel metal3 s 40542 111490 40842 111618 0 FreeSans 320 0 0 0 gpio7_6_pad_a_esd_0_h
port 2373 nsew signal bidirectional
flabel metal3 s 40542 110058 40842 110188 0 FreeSans 320 0 0 0 gpio7_6_pad_a_esd_1_h
port 2374 nsew signal bidirectional
flabel metal3 s 40542 108964 40842 109178 0 FreeSans 320 0 0 0 gpio7_6_pad_a_noesd_h
port 2375 nsew signal bidirectional
flabel metal3 s 40542 108332 40842 108402 0 FreeSans 320 0 0 0 gpio7_6_analog_en
port 2376 nsew signal input
flabel metal3 s 40542 105572 40842 105642 0 FreeSans 320 0 0 0 gpio7_6_analog_pol
port 2377 nsew signal input
flabel metal3 s 40542 104992 40842 105062 0 FreeSans 320 0 0 0 gpio7_6_inp_dis
port 2378 nsew signal input
flabel metal3 s 40542 103826 40842 103896 0 FreeSans 320 0 0 0 gpio7_6_enable_inp_h
port 2379 nsew signal input
flabel metal3 s 40542 103370 40842 103440 0 FreeSans 320 0 0 0 gpio7_6_enable_h
port 2380 nsew signal input
flabel metal3 s 40542 102916 40842 102986 0 FreeSans 320 0 0 0 gpio7_6_hld_h_n
port 2381 nsew signal input
flabel metal3 s 40542 102298 40842 102368 0 FreeSans 320 0 0 0 gpio7_6_analog_sel
port 2382 nsew signal input
flabel metal3 s 40542 101854 40842 101924 0 FreeSans 320 0 0 0 gpio7_6_dm[2]
port 2383 nsew signal input
flabel metal3 s 40542 109528 40842 109598 0 FreeSans 320 0 0 0 gpio7_6_dm[1]
port 2384 nsew signal input
flabel metal3 s 40542 106120 40842 106190 0 FreeSans 320 0 0 0 gpio7_6_dm[0]
port 2385 nsew signal input
flabel metal3 s 40542 101370 40842 101440 0 FreeSans 320 0 0 0 gpio7_6_hld_ovr
port 2386 nsew signal input
flabel metal3 s 40542 100598 40842 100668 0 FreeSans 320 0 0 0 gpio7_6_out
port 2387 nsew signal input
flabel metal3 s 40542 99398 40842 99468 0 FreeSans 320 0 0 0 gpio7_6_enable_vswitch_h
port 2388 nsew signal input
flabel metal3 s 40542 98678 40842 98748 0 FreeSans 320 0 0 0 gpio7_6_enable_vdda_h
port 2389 nsew signal input
flabel metal3 s 40542 97816 40842 97886 0 FreeSans 320 0 0 0 gpio7_6_vtrip_sel
port 2390 nsew signal input
flabel metal3 s 40542 97472 40842 97542 0 FreeSans 320 0 0 0 gpio7_6_ib_mode_sel
port 2391 nsew signal input
flabel metal3 s 40542 97062 40842 97132 0 FreeSans 320 0 0 0 gpio7_6_oe_n
port 2392 nsew signal input
flabel metal3 s 40542 96480 40842 96604 0 FreeSans 320 0 0 0 gpio7_6_in_h
port 2393 nsew signal output
flabel metal3 s 40542 114202 40842 114272 0 FreeSans 320 0 0 0 gpio7_6_zero
port 2394 nsew signal output
flabel metal3 s 40542 114652 40842 114722 0 FreeSans 320 0 0 0 gpio7_6_one
port 2395 nsew signal output
flabel metal3 s 40542 92002 40842 92072 0 FreeSans 320 0 0 0 gpio7_7_tie_lo_esd
port 2396 nsew signal output
flabel metal3 s 40538 91424 40838 91494 0 FreeSans 320 0 0 0 gpio7_7_in
port 2397 nsew signal output
flabel metal3 s 40542 91704 40842 91774 0 FreeSans 320 0 0 0 gpio7_7_tie_hi_esd
port 2398 nsew signal output
flabel metal3 s 40542 91112 40842 91182 0 FreeSans 320 0 0 0 gpio7_7_enable_vddio
port 2399 nsew signal input
flabel metal3 s 40542 90838 40842 90908 0 FreeSans 320 0 0 0 gpio7_7_slow
port 2400 nsew signal input
flabel metal3 s 40542 90490 40842 90618 0 FreeSans 320 0 0 0 gpio7_7_pad_a_esd_0_h
port 2401 nsew signal bidirectional
flabel metal3 s 40542 89058 40842 89188 0 FreeSans 320 0 0 0 gpio7_7_pad_a_esd_1_h
port 2402 nsew signal bidirectional
flabel metal3 s 40542 87964 40842 88178 0 FreeSans 320 0 0 0 gpio7_7_pad_a_noesd_h
port 2403 nsew signal bidirectional
flabel metal3 s 40542 87332 40842 87402 0 FreeSans 320 0 0 0 gpio7_7_analog_en
port 2404 nsew signal input
flabel metal3 s 40542 84572 40842 84642 0 FreeSans 320 0 0 0 gpio7_7_analog_pol
port 2405 nsew signal input
flabel metal3 s 40542 83992 40842 84062 0 FreeSans 320 0 0 0 gpio7_7_inp_dis
port 2406 nsew signal input
flabel metal3 s 40542 82826 40842 82896 0 FreeSans 320 0 0 0 gpio7_7_enable_inp_h
port 2407 nsew signal input
flabel metal3 s 40542 82370 40842 82440 0 FreeSans 320 0 0 0 gpio7_7_enable_h
port 2408 nsew signal input
flabel metal3 s 40542 81916 40842 81986 0 FreeSans 320 0 0 0 gpio7_7_hld_h_n
port 2409 nsew signal input
flabel metal3 s 40542 81298 40842 81368 0 FreeSans 320 0 0 0 gpio7_7_analog_sel
port 2410 nsew signal input
flabel metal3 s 40542 80854 40842 80924 0 FreeSans 320 0 0 0 gpio7_7_dm[2]
port 2411 nsew signal input
flabel metal3 s 40542 88528 40842 88598 0 FreeSans 320 0 0 0 gpio7_7_dm[1]
port 2412 nsew signal input
flabel metal3 s 40542 85120 40842 85190 0 FreeSans 320 0 0 0 gpio7_7_dm[0]
port 2413 nsew signal input
flabel metal3 s 40542 80370 40842 80440 0 FreeSans 320 0 0 0 gpio7_7_hld_ovr
port 2414 nsew signal input
flabel metal3 s 40542 79598 40842 79668 0 FreeSans 320 0 0 0 gpio7_7_out
port 2415 nsew signal input
flabel metal3 s 40542 78398 40842 78468 0 FreeSans 320 0 0 0 gpio7_7_enable_vswitch_h
port 2416 nsew signal input
flabel metal3 s 40542 77678 40842 77748 0 FreeSans 320 0 0 0 gpio7_7_enable_vdda_h
port 2417 nsew signal input
flabel metal3 s 40542 76816 40842 76886 0 FreeSans 320 0 0 0 gpio7_7_vtrip_sel
port 2418 nsew signal input
flabel metal3 s 40542 76472 40842 76542 0 FreeSans 320 0 0 0 gpio7_7_ib_mode_sel
port 2419 nsew signal input
flabel metal3 s 40542 76062 40842 76132 0 FreeSans 320 0 0 0 gpio7_7_oe_n
port 2420 nsew signal input
flabel metal3 s 40542 75480 40842 75604 0 FreeSans 320 0 0 0 gpio7_7_in_h
port 2421 nsew signal output
flabel metal3 s 40542 93202 40842 93272 0 FreeSans 320 0 0 0 gpio7_7_zero
port 2422 nsew signal output
flabel metal3 s 40542 93652 40842 93722 0 FreeSans 320 0 0 0 gpio7_7_one
port 2423 nsew signal output
flabel metal3 s 40600 47954 40900 48014 0 FreeSans 320 0 0 0 muxsplit_sw_hld_vdda_h_n
port 2424 nsew signal input
flabel metal3 s 40600 47074 40900 47134 0 FreeSans 320 0 0 0 muxsplit_sw_enable_vdda_h
port 2425 nsew signal input
flabel metal3 s 40600 43452 40900 43512 0 FreeSans 320 0 0 0 muxsplit_sw_switch_aa_sl
port 2426 nsew signal input
flabel metal3 s 40600 43200 40900 43260 0 FreeSans 320 0 0 0 muxsplit_sw_switch_aa_s0
port 2427 nsew signal input
flabel metal3 s 40600 42948 40900 43008 0 FreeSans 320 0 0 0 muxsplit_sw_switch_bb_s0
port 2428 nsew signal input
flabel metal3 s 40600 42696 40900 42756 0 FreeSans 320 0 0 0 muxsplit_sw_switch_bb_sl
port 2429 nsew signal input
flabel metal3 s 40600 42444 40900 42504 0 FreeSans 320 0 0 0 muxsplit_sw_switch_bb_sr
port 2430 nsew signal input
flabel metal3 s 40600 42108 40900 42168 0 FreeSans 320 0 0 0 muxsplit_sw_switch_aa_sr
port 2431 nsew signal input
flabel metal3 s 39793 954200 40793 958851 0 FreeSans 8000 90 0 0 vccd2[2]
port 158 nsew power bidirectional
<< end >>
